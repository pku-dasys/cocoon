module Dispatch(
  input  [175:0] io_configuration,
  output [10:0]  io_outs_15,
  output [10:0]  io_outs_14,
  output [10:0]  io_outs_13,
  output [10:0]  io_outs_12,
  output [10:0]  io_outs_11,
  output [10:0]  io_outs_10,
  output [10:0]  io_outs_9,
  output [10:0]  io_outs_8,
  output [10:0]  io_outs_7,
  output [10:0]  io_outs_6,
  output [10:0]  io_outs_5,
  output [10:0]  io_outs_4,
  output [10:0]  io_outs_3,
  output [10:0]  io_outs_2,
  output [10:0]  io_outs_1,
  output [10:0]  io_outs_0
);
  assign io_outs_15 = io_configuration[175:165]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_14 = io_configuration[164:154]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_13 = io_configuration[153:143]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_12 = io_configuration[142:132]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_11 = io_configuration[131:121]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_10 = io_configuration[120:110]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_9 = io_configuration[109:99]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_8 = io_configuration[98:88]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_7 = io_configuration[87:77]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_6 = io_configuration[76:66]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_5 = io_configuration[65:55]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_4 = io_configuration[54:44]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_3 = io_configuration[43:33]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_2 = io_configuration[32:22]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[21:11]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[10:0]; // @[BasicChiselModules.scala 464:18]
endmodule
module RegNextN(
  input         clock,
  input         reset,
  input  [4:0]  io_latency,
  input  [31:0] io_input,
  output [31:0] io_out
);
  reg [31:0] regArray_0; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_0;
  reg [31:0] regArray_1; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_1;
  reg [31:0] regArray_2; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_2;
  reg [31:0] regArray_3; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_3;
  reg [31:0] regArray_4; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_4;
  reg [31:0] regArray_5; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_5;
  reg [31:0] regArray_6; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_6;
  reg [31:0] regArray_7; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_7;
  reg [31:0] regArray_8; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_8;
  reg [31:0] regArray_9; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_9;
  reg [31:0] regArray_10; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_10;
  reg [31:0] regArray_11; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_11;
  reg [31:0] regArray_12; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_12;
  reg [31:0] regArray_13; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_13;
  reg [31:0] regArray_14; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_14;
  reg [31:0] regArray_15; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_15;
  reg [31:0] regArray_16; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_16;
  reg [31:0] regArray_17; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_17;
  reg [31:0] regArray_18; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_18;
  reg [31:0] regArray_19; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_19;
  reg [31:0] regArray_20; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_20;
  reg [31:0] regArray_21; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_21;
  reg [31:0] regArray_22; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_22;
  reg [31:0] regArray_23; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_23;
  reg [31:0] regArray_24; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_24;
  reg [31:0] regArray_25; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_25;
  reg [31:0] regArray_26; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_26;
  reg [31:0] regArray_27; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_27;
  reg [31:0] regArray_28; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_28;
  reg [31:0] regArray_29; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_29;
  reg [31:0] regArray_30; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_30;
  reg [31:0] regArray_31; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_31;
  reg [4:0] posReg; // @[BasicChiselModules.scala 41:23]
  reg [31:0] _RAND_32;
  wire  _T_1; // @[BasicChiselModules.scala 43:19]
  wire [4:0] _T_3; // @[BasicChiselModules.scala 44:31]
  wire [31:0] _GEN_1; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_2; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_3; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_4; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_5; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_6; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_7; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_8; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_9; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_10; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_11; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_12; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_13; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_14; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_15; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_16; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_17; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_18; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_19; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_20; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_21; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_22; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_23; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_24; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_25; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_26; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_27; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_28; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_29; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_30; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_31; // @[BasicChiselModules.scala 44:12]
  wire [4:0] _T_5; // @[BasicChiselModules.scala 49:20]
  assign _T_1 = io_latency > 5'h0; // @[BasicChiselModules.scala 43:19]
  assign _T_3 = posReg - io_latency; // @[BasicChiselModules.scala 44:31]
  assign _GEN_1 = 5'h1 == _T_3 ? regArray_1 : regArray_0; // @[BasicChiselModules.scala 44:12]
  assign _GEN_2 = 5'h2 == _T_3 ? regArray_2 : _GEN_1; // @[BasicChiselModules.scala 44:12]
  assign _GEN_3 = 5'h3 == _T_3 ? regArray_3 : _GEN_2; // @[BasicChiselModules.scala 44:12]
  assign _GEN_4 = 5'h4 == _T_3 ? regArray_4 : _GEN_3; // @[BasicChiselModules.scala 44:12]
  assign _GEN_5 = 5'h5 == _T_3 ? regArray_5 : _GEN_4; // @[BasicChiselModules.scala 44:12]
  assign _GEN_6 = 5'h6 == _T_3 ? regArray_6 : _GEN_5; // @[BasicChiselModules.scala 44:12]
  assign _GEN_7 = 5'h7 == _T_3 ? regArray_7 : _GEN_6; // @[BasicChiselModules.scala 44:12]
  assign _GEN_8 = 5'h8 == _T_3 ? regArray_8 : _GEN_7; // @[BasicChiselModules.scala 44:12]
  assign _GEN_9 = 5'h9 == _T_3 ? regArray_9 : _GEN_8; // @[BasicChiselModules.scala 44:12]
  assign _GEN_10 = 5'ha == _T_3 ? regArray_10 : _GEN_9; // @[BasicChiselModules.scala 44:12]
  assign _GEN_11 = 5'hb == _T_3 ? regArray_11 : _GEN_10; // @[BasicChiselModules.scala 44:12]
  assign _GEN_12 = 5'hc == _T_3 ? regArray_12 : _GEN_11; // @[BasicChiselModules.scala 44:12]
  assign _GEN_13 = 5'hd == _T_3 ? regArray_13 : _GEN_12; // @[BasicChiselModules.scala 44:12]
  assign _GEN_14 = 5'he == _T_3 ? regArray_14 : _GEN_13; // @[BasicChiselModules.scala 44:12]
  assign _GEN_15 = 5'hf == _T_3 ? regArray_15 : _GEN_14; // @[BasicChiselModules.scala 44:12]
  assign _GEN_16 = 5'h10 == _T_3 ? regArray_16 : _GEN_15; // @[BasicChiselModules.scala 44:12]
  assign _GEN_17 = 5'h11 == _T_3 ? regArray_17 : _GEN_16; // @[BasicChiselModules.scala 44:12]
  assign _GEN_18 = 5'h12 == _T_3 ? regArray_18 : _GEN_17; // @[BasicChiselModules.scala 44:12]
  assign _GEN_19 = 5'h13 == _T_3 ? regArray_19 : _GEN_18; // @[BasicChiselModules.scala 44:12]
  assign _GEN_20 = 5'h14 == _T_3 ? regArray_20 : _GEN_19; // @[BasicChiselModules.scala 44:12]
  assign _GEN_21 = 5'h15 == _T_3 ? regArray_21 : _GEN_20; // @[BasicChiselModules.scala 44:12]
  assign _GEN_22 = 5'h16 == _T_3 ? regArray_22 : _GEN_21; // @[BasicChiselModules.scala 44:12]
  assign _GEN_23 = 5'h17 == _T_3 ? regArray_23 : _GEN_22; // @[BasicChiselModules.scala 44:12]
  assign _GEN_24 = 5'h18 == _T_3 ? regArray_24 : _GEN_23; // @[BasicChiselModules.scala 44:12]
  assign _GEN_25 = 5'h19 == _T_3 ? regArray_25 : _GEN_24; // @[BasicChiselModules.scala 44:12]
  assign _GEN_26 = 5'h1a == _T_3 ? regArray_26 : _GEN_25; // @[BasicChiselModules.scala 44:12]
  assign _GEN_27 = 5'h1b == _T_3 ? regArray_27 : _GEN_26; // @[BasicChiselModules.scala 44:12]
  assign _GEN_28 = 5'h1c == _T_3 ? regArray_28 : _GEN_27; // @[BasicChiselModules.scala 44:12]
  assign _GEN_29 = 5'h1d == _T_3 ? regArray_29 : _GEN_28; // @[BasicChiselModules.scala 44:12]
  assign _GEN_30 = 5'h1e == _T_3 ? regArray_30 : _GEN_29; // @[BasicChiselModules.scala 44:12]
  assign _GEN_31 = 5'h1f == _T_3 ? regArray_31 : _GEN_30; // @[BasicChiselModules.scala 44:12]
  assign _T_5 = posReg + 5'h1; // @[BasicChiselModules.scala 49:20]
  assign io_out = _T_1 ? _GEN_31 : io_input; // @[BasicChiselModules.scala 44:12 BasicChiselModules.scala 47:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regArray_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regArray_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regArray_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regArray_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regArray_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regArray_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regArray_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regArray_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regArray_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regArray_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regArray_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regArray_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regArray_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regArray_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regArray_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regArray_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regArray_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regArray_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regArray_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regArray_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regArray_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regArray_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regArray_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regArray_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regArray_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regArray_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regArray_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regArray_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regArray_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regArray_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regArray_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regArray_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  posReg = _RAND_32[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regArray_0 <= 32'h0;
    end else if (_T_1) begin
      if (5'h0 == posReg) begin
        regArray_0 <= io_input;
      end
    end
    if (reset) begin
      regArray_1 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1 == posReg) begin
        regArray_1 <= io_input;
      end
    end
    if (reset) begin
      regArray_2 <= 32'h0;
    end else if (_T_1) begin
      if (5'h2 == posReg) begin
        regArray_2 <= io_input;
      end
    end
    if (reset) begin
      regArray_3 <= 32'h0;
    end else if (_T_1) begin
      if (5'h3 == posReg) begin
        regArray_3 <= io_input;
      end
    end
    if (reset) begin
      regArray_4 <= 32'h0;
    end else if (_T_1) begin
      if (5'h4 == posReg) begin
        regArray_4 <= io_input;
      end
    end
    if (reset) begin
      regArray_5 <= 32'h0;
    end else if (_T_1) begin
      if (5'h5 == posReg) begin
        regArray_5 <= io_input;
      end
    end
    if (reset) begin
      regArray_6 <= 32'h0;
    end else if (_T_1) begin
      if (5'h6 == posReg) begin
        regArray_6 <= io_input;
      end
    end
    if (reset) begin
      regArray_7 <= 32'h0;
    end else if (_T_1) begin
      if (5'h7 == posReg) begin
        regArray_7 <= io_input;
      end
    end
    if (reset) begin
      regArray_8 <= 32'h0;
    end else if (_T_1) begin
      if (5'h8 == posReg) begin
        regArray_8 <= io_input;
      end
    end
    if (reset) begin
      regArray_9 <= 32'h0;
    end else if (_T_1) begin
      if (5'h9 == posReg) begin
        regArray_9 <= io_input;
      end
    end
    if (reset) begin
      regArray_10 <= 32'h0;
    end else if (_T_1) begin
      if (5'ha == posReg) begin
        regArray_10 <= io_input;
      end
    end
    if (reset) begin
      regArray_11 <= 32'h0;
    end else if (_T_1) begin
      if (5'hb == posReg) begin
        regArray_11 <= io_input;
      end
    end
    if (reset) begin
      regArray_12 <= 32'h0;
    end else if (_T_1) begin
      if (5'hc == posReg) begin
        regArray_12 <= io_input;
      end
    end
    if (reset) begin
      regArray_13 <= 32'h0;
    end else if (_T_1) begin
      if (5'hd == posReg) begin
        regArray_13 <= io_input;
      end
    end
    if (reset) begin
      regArray_14 <= 32'h0;
    end else if (_T_1) begin
      if (5'he == posReg) begin
        regArray_14 <= io_input;
      end
    end
    if (reset) begin
      regArray_15 <= 32'h0;
    end else if (_T_1) begin
      if (5'hf == posReg) begin
        regArray_15 <= io_input;
      end
    end
    if (reset) begin
      regArray_16 <= 32'h0;
    end else if (_T_1) begin
      if (5'h10 == posReg) begin
        regArray_16 <= io_input;
      end
    end
    if (reset) begin
      regArray_17 <= 32'h0;
    end else if (_T_1) begin
      if (5'h11 == posReg) begin
        regArray_17 <= io_input;
      end
    end
    if (reset) begin
      regArray_18 <= 32'h0;
    end else if (_T_1) begin
      if (5'h12 == posReg) begin
        regArray_18 <= io_input;
      end
    end
    if (reset) begin
      regArray_19 <= 32'h0;
    end else if (_T_1) begin
      if (5'h13 == posReg) begin
        regArray_19 <= io_input;
      end
    end
    if (reset) begin
      regArray_20 <= 32'h0;
    end else if (_T_1) begin
      if (5'h14 == posReg) begin
        regArray_20 <= io_input;
      end
    end
    if (reset) begin
      regArray_21 <= 32'h0;
    end else if (_T_1) begin
      if (5'h15 == posReg) begin
        regArray_21 <= io_input;
      end
    end
    if (reset) begin
      regArray_22 <= 32'h0;
    end else if (_T_1) begin
      if (5'h16 == posReg) begin
        regArray_22 <= io_input;
      end
    end
    if (reset) begin
      regArray_23 <= 32'h0;
    end else if (_T_1) begin
      if (5'h17 == posReg) begin
        regArray_23 <= io_input;
      end
    end
    if (reset) begin
      regArray_24 <= 32'h0;
    end else if (_T_1) begin
      if (5'h18 == posReg) begin
        regArray_24 <= io_input;
      end
    end
    if (reset) begin
      regArray_25 <= 32'h0;
    end else if (_T_1) begin
      if (5'h19 == posReg) begin
        regArray_25 <= io_input;
      end
    end
    if (reset) begin
      regArray_26 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1a == posReg) begin
        regArray_26 <= io_input;
      end
    end
    if (reset) begin
      regArray_27 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1b == posReg) begin
        regArray_27 <= io_input;
      end
    end
    if (reset) begin
      regArray_28 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1c == posReg) begin
        regArray_28 <= io_input;
      end
    end
    if (reset) begin
      regArray_29 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1d == posReg) begin
        regArray_29 <= io_input;
      end
    end
    if (reset) begin
      regArray_30 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1e == posReg) begin
        regArray_30 <= io_input;
      end
    end
    if (reset) begin
      regArray_31 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1f == posReg) begin
        regArray_31 <= io_input;
      end
    end
    if (reset) begin
      posReg <= 5'h0;
    end else begin
      posReg <= _T_5;
    end
  end
endmodule
module Synchronizer(
  input         clock,
  input         reset,
  input  [5:0]  io_skewing,
  input  [31:0] io_input0,
  input  [31:0] io_input1,
  output [31:0] io_skewedInput0,
  output [31:0] io_skewedInput1
);
  wire  regNextN_clock; // @[BasicChiselModules.scala 66:24]
  wire  regNextN_reset; // @[BasicChiselModules.scala 66:24]
  wire [4:0] regNextN_io_latency; // @[BasicChiselModules.scala 66:24]
  wire [31:0] regNextN_io_input; // @[BasicChiselModules.scala 66:24]
  wire [31:0] regNextN_io_out; // @[BasicChiselModules.scala 66:24]
  wire  signal; // @[BasicChiselModules.scala 68:26]
  RegNextN regNextN ( // @[BasicChiselModules.scala 66:24]
    .clock(regNextN_clock),
    .reset(regNextN_reset),
    .io_latency(regNextN_io_latency),
    .io_input(regNextN_io_input),
    .io_out(regNextN_io_out)
  );
  assign signal = io_skewing[5]; // @[BasicChiselModules.scala 68:26]
  assign io_skewedInput0 = signal ? regNextN_io_out : io_input0; // @[BasicChiselModules.scala 73:21 BasicChiselModules.scala 78:21]
  assign io_skewedInput1 = signal ? io_input1 : regNextN_io_out; // @[BasicChiselModules.scala 74:21 BasicChiselModules.scala 77:21]
  assign regNextN_clock = clock;
  assign regNextN_reset = reset;
  assign regNextN_io_latency = io_skewing[4:0]; // @[BasicChiselModules.scala 69:23]
  assign regNextN_io_input = signal ? io_input0 : io_input1; // @[BasicChiselModules.scala 72:23 BasicChiselModules.scala 76:23]
endmodule
module Alu(
  input         clock,
  input         reset,
  input         io_en,
  input  [5:0]  io_skewing,
  input  [3:0]  io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  synchronizer_clock; // @[BasicChiselModules.scala 242:28]
  wire  synchronizer_reset; // @[BasicChiselModules.scala 242:28]
  wire [5:0] synchronizer_io_skewing; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_input0; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_input1; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_skewedInput0; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 242:28]
  wire [31:0] _T_1; // @[BasicChiselModules.scala 220:55]
  wire [31:0] _T_3; // @[BasicChiselModules.scala 221:55]
  wire [31:0] _T_4; // @[BasicChiselModules.scala 222:55]
  wire [31:0] _T_5; // @[BasicChiselModules.scala 223:54]
  wire [31:0] _T_6; // @[BasicChiselModules.scala 224:55]
  wire [63:0] _T_7; // @[BasicChiselModules.scala 225:55]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  wire [31:0] _T_11; // @[Mux.scala 68:16]
  wire  _T_12; // @[Mux.scala 68:19]
  wire [63:0] _T_13; // @[Mux.scala 68:16]
  wire  _T_14; // @[Mux.scala 68:19]
  wire [63:0] _T_15; // @[Mux.scala 68:16]
  wire  _T_16; // @[Mux.scala 68:19]
  wire [63:0] _T_17; // @[Mux.scala 68:16]
  wire  _T_18; // @[Mux.scala 68:19]
  wire [63:0] _T_19; // @[Mux.scala 68:16]
  wire  _T_20; // @[Mux.scala 68:19]
  wire [63:0] _T_21; // @[Mux.scala 68:16]
  wire  _T_22; // @[Mux.scala 68:19]
  wire [63:0] _T_23; // @[Mux.scala 68:16]
  wire [63:0] _GEN_0; // @[BasicChiselModules.scala 255:15]
  Synchronizer synchronizer ( // @[BasicChiselModules.scala 242:28]
    .clock(synchronizer_clock),
    .reset(synchronizer_reset),
    .io_skewing(synchronizer_io_skewing),
    .io_input0(synchronizer_io_input0),
    .io_input1(synchronizer_io_input1),
    .io_skewedInput0(synchronizer_io_skewedInput0),
    .io_skewedInput1(synchronizer_io_skewedInput1)
  );
  assign _T_1 = synchronizer_io_skewedInput0 + synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 220:55]
  assign _T_3 = synchronizer_io_skewedInput0 - synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 221:55]
  assign _T_4 = synchronizer_io_skewedInput0 & synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 222:55]
  assign _T_5 = synchronizer_io_skewedInput0 | synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 223:54]
  assign _T_6 = synchronizer_io_skewedInput0 ^ synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 224:55]
  assign _T_7 = synchronizer_io_skewedInput0 * synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 225:55]
  assign _T_9 = synchronizer_io_skewedInput1; // @[Mux.scala 68:16]
  assign _T_10 = 4'hc == io_configuration; // @[Mux.scala 68:19]
  assign _T_11 = _T_10 ? synchronizer_io_skewedInput0 : _T_9; // @[Mux.scala 68:16]
  assign _T_12 = 4'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_13 = _T_12 ? _T_7 : {{32'd0}, _T_11}; // @[Mux.scala 68:16]
  assign _T_14 = 4'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_15 = _T_14 ? {{32'd0}, _T_6} : _T_13; // @[Mux.scala 68:16]
  assign _T_16 = 4'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_17 = _T_16 ? {{32'd0}, _T_5} : _T_15; // @[Mux.scala 68:16]
  assign _T_18 = 4'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_19 = _T_18 ? {{32'd0}, _T_4} : _T_17; // @[Mux.scala 68:16]
  assign _T_20 = 4'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_21 = _T_20 ? {{32'd0}, _T_3} : _T_19; // @[Mux.scala 68:16]
  assign _T_22 = 4'h0 == io_configuration; // @[Mux.scala 68:19]
  assign _T_23 = _T_22 ? {{32'd0}, _T_1} : _T_21; // @[Mux.scala 68:16]
  assign _GEN_0 = io_en ? _T_23 : 64'h0; // @[BasicChiselModules.scala 255:15]
  assign io_outs_0 = _GEN_0[31:0]; // @[BasicChiselModules.scala 256:9 BasicChiselModules.scala 259:11]
  assign synchronizer_clock = clock;
  assign synchronizer_reset = reset;
  assign synchronizer_io_skewing = io_skewing; // @[BasicChiselModules.scala 246:27]
  assign synchronizer_io_input0 = io_inputs_0; // @[BasicChiselModules.scala 243:26]
  assign synchronizer_io_input1 = io_inputs_1; // @[BasicChiselModules.scala 244:26]
endmodule
module ScheduleController(
  input        clock,
  input        reset,
  input        io_en,
  input  [4:0] io_waitCycle,
  output       io_valid
);
  reg  state; // @[BasicChiselModules.scala 139:22]
  reg [31:0] _RAND_0;
  reg [4:0] cycleReg; // @[BasicChiselModules.scala 140:21]
  reg [31:0] _RAND_1;
  wire  _T; // @[BasicChiselModules.scala 142:25]
  wire  _T_2; // @[BasicChiselModules.scala 145:16]
  wire [4:0] _T_5; // @[BasicChiselModules.scala 149:30]
  wire  _GEN_0; // @[BasicChiselModules.scala 146:39]
  wire  _GEN_2; // @[BasicChiselModules.scala 145:28]
  wire  _GEN_4; // @[BasicChiselModules.scala 144:15]
  assign _T = cycleReg == io_waitCycle; // @[BasicChiselModules.scala 142:25]
  assign _T_2 = state == 1'h0; // @[BasicChiselModules.scala 145:16]
  assign _T_5 = cycleReg + 5'h1; // @[BasicChiselModules.scala 149:30]
  assign _GEN_0 = _T | state; // @[BasicChiselModules.scala 146:39]
  assign _GEN_2 = _T_2 ? _GEN_0 : state; // @[BasicChiselModules.scala 145:28]
  assign _GEN_4 = io_en & _GEN_2; // @[BasicChiselModules.scala 144:15]
  assign io_valid = _T & io_en; // @[BasicChiselModules.scala 142:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_4;
    end
    if (io_en) begin
      if (_T_2) begin
        if (!(_T)) begin
          cycleReg <= _T_5;
        end
      end
    end else begin
      cycleReg <= 5'h0;
    end
  end
endmodule
module MultiIIScheduleController(
  input         clock,
  input         reset,
  input         io_en,
  input  [10:0] io_schedules_0,
  input  [10:0] io_schedules_1,
  input  [10:0] io_schedules_2,
  input  [10:0] io_schedules_3,
  input  [1:0]  io_II,
  output        io_valid,
  output [5:0]  io_skewing
);
  wire  ScheduleController_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_io_valid; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_1_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_io_valid; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_2_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_io_valid; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_3_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_io_valid; // @[BasicChiselModules.scala 170:77]
  reg  validRegs_0; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_0;
  reg  validRegs_1; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_1;
  reg  validRegs_2; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_2;
  reg  validRegs_3; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_3;
  reg [1:0] cycleReg; // @[BasicChiselModules.scala 172:25]
  reg [31:0] _RAND_4;
  wire  _GEN_1; // @[BasicChiselModules.scala 181:12]
  wire  _GEN_2; // @[BasicChiselModules.scala 181:12]
  wire [10:0] _GEN_5; // @[BasicChiselModules.scala 182:39]
  wire [10:0] _GEN_6; // @[BasicChiselModules.scala 182:39]
  wire [10:0] _GEN_7; // @[BasicChiselModules.scala 182:39]
  wire [1:0] _T_8; // @[BasicChiselModules.scala 185:29]
  wire  _T_9; // @[BasicChiselModules.scala 185:19]
  wire [1:0] _T_11; // @[BasicChiselModules.scala 188:28]
  ScheduleController ScheduleController ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_clock),
    .reset(ScheduleController_reset),
    .io_en(ScheduleController_io_en),
    .io_waitCycle(ScheduleController_io_waitCycle),
    .io_valid(ScheduleController_io_valid)
  );
  ScheduleController ScheduleController_1 ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_1_clock),
    .reset(ScheduleController_1_reset),
    .io_en(ScheduleController_1_io_en),
    .io_waitCycle(ScheduleController_1_io_waitCycle),
    .io_valid(ScheduleController_1_io_valid)
  );
  ScheduleController ScheduleController_2 ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_2_clock),
    .reset(ScheduleController_2_reset),
    .io_en(ScheduleController_2_io_en),
    .io_waitCycle(ScheduleController_2_io_waitCycle),
    .io_valid(ScheduleController_2_io_valid)
  );
  ScheduleController ScheduleController_3 ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_3_clock),
    .reset(ScheduleController_3_reset),
    .io_en(ScheduleController_3_io_en),
    .io_waitCycle(ScheduleController_3_io_waitCycle),
    .io_valid(ScheduleController_3_io_valid)
  );
  assign _GEN_1 = 2'h1 == cycleReg ? validRegs_1 : validRegs_0; // @[BasicChiselModules.scala 181:12]
  assign _GEN_2 = 2'h2 == cycleReg ? validRegs_2 : _GEN_1; // @[BasicChiselModules.scala 181:12]
  assign _GEN_5 = 2'h1 == cycleReg ? io_schedules_1 : io_schedules_0; // @[BasicChiselModules.scala 182:39]
  assign _GEN_6 = 2'h2 == cycleReg ? io_schedules_2 : _GEN_5; // @[BasicChiselModules.scala 182:39]
  assign _GEN_7 = 2'h3 == cycleReg ? io_schedules_3 : _GEN_6; // @[BasicChiselModules.scala 182:39]
  assign _T_8 = io_II - 2'h1; // @[BasicChiselModules.scala 185:29]
  assign _T_9 = cycleReg == _T_8; // @[BasicChiselModules.scala 185:19]
  assign _T_11 = cycleReg + 2'h1; // @[BasicChiselModules.scala 188:28]
  assign io_valid = 2'h3 == cycleReg ? validRegs_3 : _GEN_2; // @[BasicChiselModules.scala 181:12]
  assign io_skewing = _GEN_7[10:5]; // @[BasicChiselModules.scala 182:14]
  assign ScheduleController_clock = clock;
  assign ScheduleController_reset = reset;
  assign ScheduleController_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_io_waitCycle = io_schedules_0[4:0]; // @[BasicChiselModules.scala 177:37]
  assign ScheduleController_1_clock = clock;
  assign ScheduleController_1_reset = reset;
  assign ScheduleController_1_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_1_io_waitCycle = io_schedules_1[4:0]; // @[BasicChiselModules.scala 177:37]
  assign ScheduleController_2_clock = clock;
  assign ScheduleController_2_reset = reset;
  assign ScheduleController_2_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_2_io_waitCycle = io_schedules_2[4:0]; // @[BasicChiselModules.scala 177:37]
  assign ScheduleController_3_clock = clock;
  assign ScheduleController_3_reset = reset;
  assign ScheduleController_3_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_3_io_waitCycle = io_schedules_3[4:0]; // @[BasicChiselModules.scala 177:37]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validRegs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  validRegs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  validRegs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  validRegs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cycleReg = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      validRegs_0 <= 1'h0;
    end else begin
      validRegs_0 <= ScheduleController_io_valid;
    end
    if (reset) begin
      validRegs_1 <= 1'h0;
    end else begin
      validRegs_1 <= ScheduleController_1_io_valid;
    end
    if (reset) begin
      validRegs_2 <= 1'h0;
    end else begin
      validRegs_2 <= ScheduleController_2_io_valid;
    end
    if (reset) begin
      validRegs_3 <= 1'h0;
    end else begin
      validRegs_3 <= ScheduleController_3_io_valid;
    end
    if (reset) begin
      cycleReg <= 2'h3;
    end else if (io_en) begin
      if (_T_9) begin
        cycleReg <= 2'h0;
      end else begin
        cycleReg <= _T_11;
      end
    end
  end
endmodule
module Dispatch_1(
  input  [2:0] io_configuration,
  output       io_outs_2,
  output       io_outs_1,
  output       io_outs_0
);
  assign io_outs_2 = io_configuration[2]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[1]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[0]; // @[BasicChiselModules.scala 464:18]
endmodule
module RegisterFile(
  input         clock,
  input         reset,
  input  [3:0]  io_configuration,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_1,
  output [31:0] io_outs_0
);
  wire [2:0] Dispatch_io_configuration; // @[BasicChiselModules.scala 332:26]
  wire  Dispatch_io_outs_2; // @[BasicChiselModules.scala 332:26]
  wire  Dispatch_io_outs_1; // @[BasicChiselModules.scala 332:26]
  wire  Dispatch_io_outs_0; // @[BasicChiselModules.scala 332:26]
  wire  _T_1; // @[BasicChiselModules.scala 336:37]
  reg [31:0] _T_3_0; // @[BasicChiselModules.scala 338:23]
  reg [31:0] _RAND_0;
  reg [31:0] _T_3_1; // @[BasicChiselModules.scala 338:23]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[BasicChiselModules.scala 340:20]
  Dispatch_1 Dispatch ( // @[BasicChiselModules.scala 332:26]
    .io_configuration(Dispatch_io_configuration),
    .io_outs_2(Dispatch_io_outs_2),
    .io_outs_1(Dispatch_io_outs_1),
    .io_outs_0(Dispatch_io_outs_0)
  );
  assign _T_1 = io_configuration[3]; // @[BasicChiselModules.scala 336:37]
  assign _T_4 = _T_1 == 1'h0; // @[BasicChiselModules.scala 340:20]
  assign io_outs_1 = Dispatch_io_outs_2 ? _T_3_1 : _T_3_0; // @[BasicChiselModules.scala 346:18]
  assign io_outs_0 = Dispatch_io_outs_1 ? _T_3_1 : _T_3_0; // @[BasicChiselModules.scala 346:18]
  assign Dispatch_io_configuration = io_configuration[2:0]; // @[BasicChiselModules.scala 334:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3_0 <= 32'h0;
    end else if (_T_4) begin
      if (1'h0 == Dispatch_io_outs_0) begin
        _T_3_0 <= io_inputs_0;
      end
    end
    if (reset) begin
      _T_3_1 <= 32'h0;
    end else if (_T_4) begin
      if (Dispatch_io_outs_0) begin
        _T_3_1 <= io_inputs_0;
      end
    end
  end
endmodule
module Multiplexer(
  input         io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  assign _T_1 = io_configuration ? io_inputs_1 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 1'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_2 ? io_inputs_0 : _T_1; // @[BasicChiselModules.scala 370:14]
endmodule
module Multiplexer_3(
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_5,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  assign _T = 3'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_5 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_4 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_3 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_2 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_9 = _T_8 ? io_inputs_1 : _T_7; // @[Mux.scala 68:16]
  assign _T_10 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_10 ? io_inputs_0 : _T_9; // @[BasicChiselModules.scala 370:14]
endmodule
module Multiplexer_4(
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  assign _T = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_4 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_3 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_1 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_8 ? io_inputs_0 : _T_7; // @[BasicChiselModules.scala 370:14]
endmodule
module Multiplexer_5(
  input  [1:0]  io_configuration,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  assign _T = 2'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_3 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 2'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_2 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 2'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_1 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 2'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_6 ? io_inputs_0 : _T_5; // @[BasicChiselModules.scala 370:14]
endmodule
module ConstUnit(
  input  [31:0] io_configuration,
  output [31:0] io_outs_0
);
  assign io_outs_0 = io_configuration; // @[BasicChiselModules.scala 403:14]
endmodule
module ConfigController(
  input        clock,
  input        reset,
  input        io_en,
  input  [1:0] io_II,
  input  [2:0] io_inConfig,
  output [2:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 96:22]
  reg [31:0] _RAND_0;
  reg [1:0] cycleReg; // @[BasicChiselModules.scala 97:21]
  reg [31:0] _RAND_1;
  reg [2:0] configRegs_0; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_2;
  reg [2:0] configRegs_1; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_3;
  reg [2:0] configRegs_2; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_4;
  reg [2:0] configRegs_3; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_5;
  wire  _T_1; // @[BasicChiselModules.scala 103:14]
  wire [2:0] _GEN_1; // @[BasicChiselModules.scala 106:18]
  wire [2:0] _GEN_2; // @[BasicChiselModules.scala 106:18]
  wire [2:0] _GEN_3; // @[BasicChiselModules.scala 106:18]
  wire  _T_3; // @[BasicChiselModules.scala 112:21]
  wire [1:0] _T_5; // @[BasicChiselModules.scala 116:30]
  wire  _GEN_9; // @[BasicChiselModules.scala 112:32]
  wire [1:0] _T_7; // @[BasicChiselModules.scala 119:31]
  wire  _T_8; // @[BasicChiselModules.scala 119:21]
  wire  _GEN_16; // @[BasicChiselModules.scala 110:34]
  wire  _GEN_22; // @[BasicChiselModules.scala 109:15]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 103:14]
  assign _GEN_1 = 2'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 106:18]
  assign _GEN_2 = 2'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 106:18]
  assign _GEN_3 = 2'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 106:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 112:21]
  assign _T_5 = cycleReg + 2'h1; // @[BasicChiselModules.scala 116:30]
  assign _GEN_9 = _T_3 | state; // @[BasicChiselModules.scala 112:32]
  assign _T_7 = io_II - 2'h1; // @[BasicChiselModules.scala 119:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 119:21]
  assign _GEN_16 = _T_1 ? _GEN_9 : state; // @[BasicChiselModules.scala 110:34]
  assign _GEN_22 = io_en & _GEN_16; // @[BasicChiselModules.scala 109:15]
  assign io_outConfig = _T_1 ? 3'h0 : _GEN_3; // @[BasicChiselModules.scala 104:18 BasicChiselModules.scala 106:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  configRegs_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  configRegs_1 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  configRegs_2 = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  configRegs_3 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_22;
    end
    if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 2'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 2'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 2'h0;
    end
    if (reset) begin
      configRegs_0 <= 3'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h0 == cycleReg) begin
          configRegs_0 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 3'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h1 == cycleReg) begin
          configRegs_1 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 3'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h2 == cycleReg) begin
          configRegs_2 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 3'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h3 == cycleReg) begin
          configRegs_3 <= io_inConfig;
        end
      end
    end
  end
endmodule
module ConfigController_1(
  input         clock,
  input         reset,
  input         io_en,
  input  [1:0]  io_II,
  input  [48:0] io_inConfig,
  output [48:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 96:22]
  reg [31:0] _RAND_0;
  reg [1:0] cycleReg; // @[BasicChiselModules.scala 97:21]
  reg [31:0] _RAND_1;
  reg [48:0] configRegs_0; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_2;
  reg [48:0] configRegs_1; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_3;
  reg [48:0] configRegs_2; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_4;
  reg [48:0] configRegs_3; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_5;
  wire  _T_1; // @[BasicChiselModules.scala 103:14]
  wire [48:0] _GEN_1; // @[BasicChiselModules.scala 106:18]
  wire [48:0] _GEN_2; // @[BasicChiselModules.scala 106:18]
  wire [48:0] _GEN_3; // @[BasicChiselModules.scala 106:18]
  wire  _T_3; // @[BasicChiselModules.scala 112:21]
  wire [1:0] _T_5; // @[BasicChiselModules.scala 116:30]
  wire  _GEN_9; // @[BasicChiselModules.scala 112:32]
  wire [1:0] _T_7; // @[BasicChiselModules.scala 119:31]
  wire  _T_8; // @[BasicChiselModules.scala 119:21]
  wire  _GEN_16; // @[BasicChiselModules.scala 110:34]
  wire  _GEN_22; // @[BasicChiselModules.scala 109:15]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 103:14]
  assign _GEN_1 = 2'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 106:18]
  assign _GEN_2 = 2'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 106:18]
  assign _GEN_3 = 2'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 106:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 112:21]
  assign _T_5 = cycleReg + 2'h1; // @[BasicChiselModules.scala 116:30]
  assign _GEN_9 = _T_3 | state; // @[BasicChiselModules.scala 112:32]
  assign _T_7 = io_II - 2'h1; // @[BasicChiselModules.scala 119:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 119:21]
  assign _GEN_16 = _T_1 ? _GEN_9 : state; // @[BasicChiselModules.scala 110:34]
  assign _GEN_22 = io_en & _GEN_16; // @[BasicChiselModules.scala 109:15]
  assign io_outConfig = _T_1 ? 49'h0 : _GEN_3; // @[BasicChiselModules.scala 104:18 BasicChiselModules.scala 106:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  configRegs_0 = _RAND_2[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  configRegs_1 = _RAND_3[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  configRegs_2 = _RAND_4[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  configRegs_3 = _RAND_5[48:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_22;
    end
    if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 2'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 2'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 2'h0;
    end
    if (reset) begin
      configRegs_0 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h0 == cycleReg) begin
          configRegs_0 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h1 == cycleReg) begin
          configRegs_1 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h2 == cycleReg) begin
          configRegs_2 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h3 == cycleReg) begin
          configRegs_3 <= io_inConfig;
        end
      end
    end
  end
endmodule
module Dispatch_6(
  input  [48:0] io_configuration,
  output [31:0] io_outs_6,
  output        io_outs_5,
  output [1:0]  io_outs_4,
  output [2:0]  io_outs_3,
  output [2:0]  io_outs_2,
  output [3:0]  io_outs_1,
  output [3:0]  io_outs_0
);
  assign io_outs_6 = io_configuration[48:17]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_5 = io_configuration[16]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_4 = io_configuration[15:14]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_3 = io_configuration[13:11]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_2 = io_configuration[10:8]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[7:4]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[3:0]; // @[BasicChiselModules.scala 464:18]
endmodule
module Dispatch_10(
  input  [198:0] io_configuration,
  output [48:0]  io_outs_4,
  output [48:0]  io_outs_3,
  output [48:0]  io_outs_2,
  output [48:0]  io_outs_1,
  output [2:0]   io_outs_0
);
  assign io_outs_4 = io_configuration[198:150]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_3 = io_configuration[149:101]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_2 = io_configuration[100:52]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[51:3]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[2:0]; // @[BasicChiselModules.scala 464:18]
endmodule
module TopModule(
  input          clock,
  input          reset,
  input          io_enConfig,
  input          io_en,
  input  [175:0] io_schedules,
  input  [1:0]   io_II,
  input  [198:0] io_configuration,
  input  [31:0]  io_inputs_1,
  input  [31:0]  io_inputs_0,
  output [31:0]  io_outs_0
);
  wire [175:0] scheduleDispatch_io_configuration; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_15; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_14; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_13; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_12; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_11; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_10; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_9; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_8; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_7; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_6; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_5; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_4; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_3; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_2; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_1; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_0; // @[TopModule.scala 119:32]
  wire  Alu_clock; // @[TopModule.scala 124:54]
  wire  Alu_reset; // @[TopModule.scala 124:54]
  wire  Alu_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_1_clock; // @[TopModule.scala 124:54]
  wire  Alu_1_reset; // @[TopModule.scala 124:54]
  wire  Alu_1_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_1_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_1_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_1_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_1_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_1_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_2_clock; // @[TopModule.scala 124:54]
  wire  Alu_2_reset; // @[TopModule.scala 124:54]
  wire  Alu_2_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_2_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_2_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_2_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_2_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_2_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_3_clock; // @[TopModule.scala 124:54]
  wire  Alu_3_reset; // @[TopModule.scala 124:54]
  wire  Alu_3_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_3_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_3_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_3_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_3_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_3_io_outs_0; // @[TopModule.scala 124:54]
  wire  MultiIIScheduleController_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_1_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_2_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_3_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 126:72]
  wire  RegisterFile_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_1_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_1_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_1_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_1_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_1_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_1_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_2_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_2_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_2_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_2_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_2_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_2_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_3_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_3_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_3_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_3_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_3_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_3_io_outs_0; // @[TopModule.scala 142:21]
  wire  Multiplexer_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_1_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_1_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_1_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_1_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_2_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_2_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_2_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_2_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_3_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_4_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_5_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_6_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_7_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_8_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_9_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_10_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_11_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_12_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_13_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_14_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_15_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_16_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_17_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_18_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_outs_0; // @[TopModule.scala 153:11]
  wire [31:0] ConstUnit_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_1_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_1_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_2_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_2_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_3_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_3_io_outs_0; // @[TopModule.scala 161:21]
  wire  configControllers_0_clock; // @[TopModule.scala 234:34]
  wire  configControllers_0_reset; // @[TopModule.scala 234:34]
  wire  configControllers_0_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_0_io_II; // @[TopModule.scala 234:34]
  wire [2:0] configControllers_0_io_inConfig; // @[TopModule.scala 234:34]
  wire [2:0] configControllers_0_io_outConfig; // @[TopModule.scala 234:34]
  wire [2:0] Dispatch_io_configuration; // @[TopModule.scala 239:26]
  wire  Dispatch_io_outs_2; // @[TopModule.scala 239:26]
  wire  Dispatch_io_outs_1; // @[TopModule.scala 239:26]
  wire  Dispatch_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_1_clock; // @[TopModule.scala 234:34]
  wire  configControllers_1_reset; // @[TopModule.scala 234:34]
  wire  configControllers_1_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_1_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_1_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_1_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_1_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_1_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_1_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_1_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_1_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_1_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_1_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_1_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_2_clock; // @[TopModule.scala 234:34]
  wire  configControllers_2_reset; // @[TopModule.scala 234:34]
  wire  configControllers_2_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_2_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_2_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_2_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_2_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_2_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_2_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_2_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_2_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_2_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_2_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_2_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_3_clock; // @[TopModule.scala 234:34]
  wire  configControllers_3_reset; // @[TopModule.scala 234:34]
  wire  configControllers_3_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_3_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_3_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_3_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_3_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_3_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_3_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_3_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_3_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_3_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_3_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_3_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_4_clock; // @[TopModule.scala 234:34]
  wire  configControllers_4_reset; // @[TopModule.scala 234:34]
  wire  configControllers_4_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_4_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_4_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_4_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_4_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_4_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_4_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_4_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_4_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_4_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_4_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_4_io_outs_0; // @[TopModule.scala 239:26]
  wire [198:0] topDispatch_io_configuration; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_4; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_3; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_2; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_1; // @[TopModule.scala 248:27]
  wire [2:0] topDispatch_io_outs_0; // @[TopModule.scala 248:27]
  Dispatch scheduleDispatch ( // @[TopModule.scala 119:32]
    .io_configuration(scheduleDispatch_io_configuration),
    .io_outs_15(scheduleDispatch_io_outs_15),
    .io_outs_14(scheduleDispatch_io_outs_14),
    .io_outs_13(scheduleDispatch_io_outs_13),
    .io_outs_12(scheduleDispatch_io_outs_12),
    .io_outs_11(scheduleDispatch_io_outs_11),
    .io_outs_10(scheduleDispatch_io_outs_10),
    .io_outs_9(scheduleDispatch_io_outs_9),
    .io_outs_8(scheduleDispatch_io_outs_8),
    .io_outs_7(scheduleDispatch_io_outs_7),
    .io_outs_6(scheduleDispatch_io_outs_6),
    .io_outs_5(scheduleDispatch_io_outs_5),
    .io_outs_4(scheduleDispatch_io_outs_4),
    .io_outs_3(scheduleDispatch_io_outs_3),
    .io_outs_2(scheduleDispatch_io_outs_2),
    .io_outs_1(scheduleDispatch_io_outs_1),
    .io_outs_0(scheduleDispatch_io_outs_0)
  );
  Alu Alu ( // @[TopModule.scala 124:54]
    .clock(Alu_clock),
    .reset(Alu_reset),
    .io_en(Alu_io_en),
    .io_skewing(Alu_io_skewing),
    .io_configuration(Alu_io_configuration),
    .io_inputs_1(Alu_io_inputs_1),
    .io_inputs_0(Alu_io_inputs_0),
    .io_outs_0(Alu_io_outs_0)
  );
  Alu Alu_1 ( // @[TopModule.scala 124:54]
    .clock(Alu_1_clock),
    .reset(Alu_1_reset),
    .io_en(Alu_1_io_en),
    .io_skewing(Alu_1_io_skewing),
    .io_configuration(Alu_1_io_configuration),
    .io_inputs_1(Alu_1_io_inputs_1),
    .io_inputs_0(Alu_1_io_inputs_0),
    .io_outs_0(Alu_1_io_outs_0)
  );
  Alu Alu_2 ( // @[TopModule.scala 124:54]
    .clock(Alu_2_clock),
    .reset(Alu_2_reset),
    .io_en(Alu_2_io_en),
    .io_skewing(Alu_2_io_skewing),
    .io_configuration(Alu_2_io_configuration),
    .io_inputs_1(Alu_2_io_inputs_1),
    .io_inputs_0(Alu_2_io_inputs_0),
    .io_outs_0(Alu_2_io_outs_0)
  );
  Alu Alu_3 ( // @[TopModule.scala 124:54]
    .clock(Alu_3_clock),
    .reset(Alu_3_reset),
    .io_en(Alu_3_io_en),
    .io_skewing(Alu_3_io_skewing),
    .io_configuration(Alu_3_io_configuration),
    .io_inputs_1(Alu_3_io_inputs_1),
    .io_inputs_0(Alu_3_io_inputs_0),
    .io_outs_0(Alu_3_io_outs_0)
  );
  MultiIIScheduleController MultiIIScheduleController ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_clock),
    .reset(MultiIIScheduleController_reset),
    .io_en(MultiIIScheduleController_io_en),
    .io_schedules_0(MultiIIScheduleController_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_io_schedules_3),
    .io_II(MultiIIScheduleController_io_II),
    .io_valid(MultiIIScheduleController_io_valid),
    .io_skewing(MultiIIScheduleController_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_1 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_1_clock),
    .reset(MultiIIScheduleController_1_reset),
    .io_en(MultiIIScheduleController_1_io_en),
    .io_schedules_0(MultiIIScheduleController_1_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_1_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_1_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_1_io_schedules_3),
    .io_II(MultiIIScheduleController_1_io_II),
    .io_valid(MultiIIScheduleController_1_io_valid),
    .io_skewing(MultiIIScheduleController_1_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_2 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_2_clock),
    .reset(MultiIIScheduleController_2_reset),
    .io_en(MultiIIScheduleController_2_io_en),
    .io_schedules_0(MultiIIScheduleController_2_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_2_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_2_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_2_io_schedules_3),
    .io_II(MultiIIScheduleController_2_io_II),
    .io_valid(MultiIIScheduleController_2_io_valid),
    .io_skewing(MultiIIScheduleController_2_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_3 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_3_clock),
    .reset(MultiIIScheduleController_3_reset),
    .io_en(MultiIIScheduleController_3_io_en),
    .io_schedules_0(MultiIIScheduleController_3_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_3_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_3_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_3_io_schedules_3),
    .io_II(MultiIIScheduleController_3_io_II),
    .io_valid(MultiIIScheduleController_3_io_valid),
    .io_skewing(MultiIIScheduleController_3_io_skewing)
  );
  RegisterFile RegisterFile ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_clock),
    .reset(RegisterFile_reset),
    .io_configuration(RegisterFile_io_configuration),
    .io_inputs_0(RegisterFile_io_inputs_0),
    .io_outs_1(RegisterFile_io_outs_1),
    .io_outs_0(RegisterFile_io_outs_0)
  );
  RegisterFile RegisterFile_1 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_1_clock),
    .reset(RegisterFile_1_reset),
    .io_configuration(RegisterFile_1_io_configuration),
    .io_inputs_0(RegisterFile_1_io_inputs_0),
    .io_outs_1(RegisterFile_1_io_outs_1),
    .io_outs_0(RegisterFile_1_io_outs_0)
  );
  RegisterFile RegisterFile_2 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_2_clock),
    .reset(RegisterFile_2_reset),
    .io_configuration(RegisterFile_2_io_configuration),
    .io_inputs_0(RegisterFile_2_io_inputs_0),
    .io_outs_1(RegisterFile_2_io_outs_1),
    .io_outs_0(RegisterFile_2_io_outs_0)
  );
  RegisterFile RegisterFile_3 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_3_clock),
    .reset(RegisterFile_3_reset),
    .io_configuration(RegisterFile_3_io_configuration),
    .io_inputs_0(RegisterFile_3_io_inputs_0),
    .io_outs_1(RegisterFile_3_io_outs_1),
    .io_outs_0(RegisterFile_3_io_outs_0)
  );
  Multiplexer Multiplexer ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_io_configuration),
    .io_inputs_1(Multiplexer_io_inputs_1),
    .io_inputs_0(Multiplexer_io_inputs_0),
    .io_outs_0(Multiplexer_io_outs_0)
  );
  Multiplexer Multiplexer_1 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_1_io_configuration),
    .io_inputs_1(Multiplexer_1_io_inputs_1),
    .io_inputs_0(Multiplexer_1_io_inputs_0),
    .io_outs_0(Multiplexer_1_io_outs_0)
  );
  Multiplexer Multiplexer_2 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_2_io_configuration),
    .io_inputs_1(Multiplexer_2_io_inputs_1),
    .io_inputs_0(Multiplexer_2_io_inputs_0),
    .io_outs_0(Multiplexer_2_io_outs_0)
  );
  Multiplexer_3 Multiplexer_3 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_3_io_configuration),
    .io_inputs_5(Multiplexer_3_io_inputs_5),
    .io_inputs_4(Multiplexer_3_io_inputs_4),
    .io_inputs_3(Multiplexer_3_io_inputs_3),
    .io_inputs_2(Multiplexer_3_io_inputs_2),
    .io_inputs_1(Multiplexer_3_io_inputs_1),
    .io_inputs_0(Multiplexer_3_io_inputs_0),
    .io_outs_0(Multiplexer_3_io_outs_0)
  );
  Multiplexer_4 Multiplexer_4 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_4_io_configuration),
    .io_inputs_4(Multiplexer_4_io_inputs_4),
    .io_inputs_3(Multiplexer_4_io_inputs_3),
    .io_inputs_2(Multiplexer_4_io_inputs_2),
    .io_inputs_1(Multiplexer_4_io_inputs_1),
    .io_inputs_0(Multiplexer_4_io_inputs_0),
    .io_outs_0(Multiplexer_4_io_outs_0)
  );
  Multiplexer_5 Multiplexer_5 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_5_io_configuration),
    .io_inputs_3(Multiplexer_5_io_inputs_3),
    .io_inputs_2(Multiplexer_5_io_inputs_2),
    .io_inputs_1(Multiplexer_5_io_inputs_1),
    .io_inputs_0(Multiplexer_5_io_inputs_0),
    .io_outs_0(Multiplexer_5_io_outs_0)
  );
  Multiplexer Multiplexer_6 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_6_io_configuration),
    .io_inputs_1(Multiplexer_6_io_inputs_1),
    .io_inputs_0(Multiplexer_6_io_inputs_0),
    .io_outs_0(Multiplexer_6_io_outs_0)
  );
  Multiplexer_3 Multiplexer_7 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_7_io_configuration),
    .io_inputs_5(Multiplexer_7_io_inputs_5),
    .io_inputs_4(Multiplexer_7_io_inputs_4),
    .io_inputs_3(Multiplexer_7_io_inputs_3),
    .io_inputs_2(Multiplexer_7_io_inputs_2),
    .io_inputs_1(Multiplexer_7_io_inputs_1),
    .io_inputs_0(Multiplexer_7_io_inputs_0),
    .io_outs_0(Multiplexer_7_io_outs_0)
  );
  Multiplexer_4 Multiplexer_8 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_8_io_configuration),
    .io_inputs_4(Multiplexer_8_io_inputs_4),
    .io_inputs_3(Multiplexer_8_io_inputs_3),
    .io_inputs_2(Multiplexer_8_io_inputs_2),
    .io_inputs_1(Multiplexer_8_io_inputs_1),
    .io_inputs_0(Multiplexer_8_io_inputs_0),
    .io_outs_0(Multiplexer_8_io_outs_0)
  );
  Multiplexer_5 Multiplexer_9 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_9_io_configuration),
    .io_inputs_3(Multiplexer_9_io_inputs_3),
    .io_inputs_2(Multiplexer_9_io_inputs_2),
    .io_inputs_1(Multiplexer_9_io_inputs_1),
    .io_inputs_0(Multiplexer_9_io_inputs_0),
    .io_outs_0(Multiplexer_9_io_outs_0)
  );
  Multiplexer Multiplexer_10 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_10_io_configuration),
    .io_inputs_1(Multiplexer_10_io_inputs_1),
    .io_inputs_0(Multiplexer_10_io_inputs_0),
    .io_outs_0(Multiplexer_10_io_outs_0)
  );
  Multiplexer_3 Multiplexer_11 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_11_io_configuration),
    .io_inputs_5(Multiplexer_11_io_inputs_5),
    .io_inputs_4(Multiplexer_11_io_inputs_4),
    .io_inputs_3(Multiplexer_11_io_inputs_3),
    .io_inputs_2(Multiplexer_11_io_inputs_2),
    .io_inputs_1(Multiplexer_11_io_inputs_1),
    .io_inputs_0(Multiplexer_11_io_inputs_0),
    .io_outs_0(Multiplexer_11_io_outs_0)
  );
  Multiplexer_4 Multiplexer_12 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_12_io_configuration),
    .io_inputs_4(Multiplexer_12_io_inputs_4),
    .io_inputs_3(Multiplexer_12_io_inputs_3),
    .io_inputs_2(Multiplexer_12_io_inputs_2),
    .io_inputs_1(Multiplexer_12_io_inputs_1),
    .io_inputs_0(Multiplexer_12_io_inputs_0),
    .io_outs_0(Multiplexer_12_io_outs_0)
  );
  Multiplexer_5 Multiplexer_13 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_13_io_configuration),
    .io_inputs_3(Multiplexer_13_io_inputs_3),
    .io_inputs_2(Multiplexer_13_io_inputs_2),
    .io_inputs_1(Multiplexer_13_io_inputs_1),
    .io_inputs_0(Multiplexer_13_io_inputs_0),
    .io_outs_0(Multiplexer_13_io_outs_0)
  );
  Multiplexer Multiplexer_14 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_14_io_configuration),
    .io_inputs_1(Multiplexer_14_io_inputs_1),
    .io_inputs_0(Multiplexer_14_io_inputs_0),
    .io_outs_0(Multiplexer_14_io_outs_0)
  );
  Multiplexer_3 Multiplexer_15 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_15_io_configuration),
    .io_inputs_5(Multiplexer_15_io_inputs_5),
    .io_inputs_4(Multiplexer_15_io_inputs_4),
    .io_inputs_3(Multiplexer_15_io_inputs_3),
    .io_inputs_2(Multiplexer_15_io_inputs_2),
    .io_inputs_1(Multiplexer_15_io_inputs_1),
    .io_inputs_0(Multiplexer_15_io_inputs_0),
    .io_outs_0(Multiplexer_15_io_outs_0)
  );
  Multiplexer_4 Multiplexer_16 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_16_io_configuration),
    .io_inputs_4(Multiplexer_16_io_inputs_4),
    .io_inputs_3(Multiplexer_16_io_inputs_3),
    .io_inputs_2(Multiplexer_16_io_inputs_2),
    .io_inputs_1(Multiplexer_16_io_inputs_1),
    .io_inputs_0(Multiplexer_16_io_inputs_0),
    .io_outs_0(Multiplexer_16_io_outs_0)
  );
  Multiplexer_5 Multiplexer_17 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_17_io_configuration),
    .io_inputs_3(Multiplexer_17_io_inputs_3),
    .io_inputs_2(Multiplexer_17_io_inputs_2),
    .io_inputs_1(Multiplexer_17_io_inputs_1),
    .io_inputs_0(Multiplexer_17_io_inputs_0),
    .io_outs_0(Multiplexer_17_io_outs_0)
  );
  Multiplexer Multiplexer_18 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_18_io_configuration),
    .io_inputs_1(Multiplexer_18_io_inputs_1),
    .io_inputs_0(Multiplexer_18_io_inputs_0),
    .io_outs_0(Multiplexer_18_io_outs_0)
  );
  ConstUnit ConstUnit ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_io_configuration),
    .io_outs_0(ConstUnit_io_outs_0)
  );
  ConstUnit ConstUnit_1 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_1_io_configuration),
    .io_outs_0(ConstUnit_1_io_outs_0)
  );
  ConstUnit ConstUnit_2 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_2_io_configuration),
    .io_outs_0(ConstUnit_2_io_outs_0)
  );
  ConstUnit ConstUnit_3 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_3_io_configuration),
    .io_outs_0(ConstUnit_3_io_outs_0)
  );
  ConfigController configControllers_0 ( // @[TopModule.scala 234:34]
    .clock(configControllers_0_clock),
    .reset(configControllers_0_reset),
    .io_en(configControllers_0_io_en),
    .io_II(configControllers_0_io_II),
    .io_inConfig(configControllers_0_io_inConfig),
    .io_outConfig(configControllers_0_io_outConfig)
  );
  Dispatch_1 Dispatch ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_io_configuration),
    .io_outs_2(Dispatch_io_outs_2),
    .io_outs_1(Dispatch_io_outs_1),
    .io_outs_0(Dispatch_io_outs_0)
  );
  ConfigController_1 configControllers_1 ( // @[TopModule.scala 234:34]
    .clock(configControllers_1_clock),
    .reset(configControllers_1_reset),
    .io_en(configControllers_1_io_en),
    .io_II(configControllers_1_io_II),
    .io_inConfig(configControllers_1_io_inConfig),
    .io_outConfig(configControllers_1_io_outConfig)
  );
  Dispatch_6 Dispatch_1 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_1_io_configuration),
    .io_outs_6(Dispatch_1_io_outs_6),
    .io_outs_5(Dispatch_1_io_outs_5),
    .io_outs_4(Dispatch_1_io_outs_4),
    .io_outs_3(Dispatch_1_io_outs_3),
    .io_outs_2(Dispatch_1_io_outs_2),
    .io_outs_1(Dispatch_1_io_outs_1),
    .io_outs_0(Dispatch_1_io_outs_0)
  );
  ConfigController_1 configControllers_2 ( // @[TopModule.scala 234:34]
    .clock(configControllers_2_clock),
    .reset(configControllers_2_reset),
    .io_en(configControllers_2_io_en),
    .io_II(configControllers_2_io_II),
    .io_inConfig(configControllers_2_io_inConfig),
    .io_outConfig(configControllers_2_io_outConfig)
  );
  Dispatch_6 Dispatch_2 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_2_io_configuration),
    .io_outs_6(Dispatch_2_io_outs_6),
    .io_outs_5(Dispatch_2_io_outs_5),
    .io_outs_4(Dispatch_2_io_outs_4),
    .io_outs_3(Dispatch_2_io_outs_3),
    .io_outs_2(Dispatch_2_io_outs_2),
    .io_outs_1(Dispatch_2_io_outs_1),
    .io_outs_0(Dispatch_2_io_outs_0)
  );
  ConfigController_1 configControllers_3 ( // @[TopModule.scala 234:34]
    .clock(configControllers_3_clock),
    .reset(configControllers_3_reset),
    .io_en(configControllers_3_io_en),
    .io_II(configControllers_3_io_II),
    .io_inConfig(configControllers_3_io_inConfig),
    .io_outConfig(configControllers_3_io_outConfig)
  );
  Dispatch_6 Dispatch_3 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_3_io_configuration),
    .io_outs_6(Dispatch_3_io_outs_6),
    .io_outs_5(Dispatch_3_io_outs_5),
    .io_outs_4(Dispatch_3_io_outs_4),
    .io_outs_3(Dispatch_3_io_outs_3),
    .io_outs_2(Dispatch_3_io_outs_2),
    .io_outs_1(Dispatch_3_io_outs_1),
    .io_outs_0(Dispatch_3_io_outs_0)
  );
  ConfigController_1 configControllers_4 ( // @[TopModule.scala 234:34]
    .clock(configControllers_4_clock),
    .reset(configControllers_4_reset),
    .io_en(configControllers_4_io_en),
    .io_II(configControllers_4_io_II),
    .io_inConfig(configControllers_4_io_inConfig),
    .io_outConfig(configControllers_4_io_outConfig)
  );
  Dispatch_6 Dispatch_4 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_4_io_configuration),
    .io_outs_6(Dispatch_4_io_outs_6),
    .io_outs_5(Dispatch_4_io_outs_5),
    .io_outs_4(Dispatch_4_io_outs_4),
    .io_outs_3(Dispatch_4_io_outs_3),
    .io_outs_2(Dispatch_4_io_outs_2),
    .io_outs_1(Dispatch_4_io_outs_1),
    .io_outs_0(Dispatch_4_io_outs_0)
  );
  Dispatch_10 topDispatch ( // @[TopModule.scala 248:27]
    .io_configuration(topDispatch_io_configuration),
    .io_outs_4(topDispatch_io_outs_4),
    .io_outs_3(topDispatch_io_outs_3),
    .io_outs_2(topDispatch_io_outs_2),
    .io_outs_1(topDispatch_io_outs_1),
    .io_outs_0(topDispatch_io_outs_0)
  );
  assign io_outs_0 = Multiplexer_io_outs_0; // @[TopModule.scala 263:25]
  assign scheduleDispatch_io_configuration = io_schedules; // @[TopModule.scala 120:37]
  assign Alu_clock = clock;
  assign Alu_reset = reset;
  assign Alu_io_en = MultiIIScheduleController_io_valid; // @[TopModule.scala 135:15]
  assign Alu_io_skewing = MultiIIScheduleController_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_io_configuration = Dispatch_1_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_io_inputs_1 = Multiplexer_4_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_io_inputs_0 = Multiplexer_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_1_clock = clock;
  assign Alu_1_reset = reset;
  assign Alu_1_io_en = MultiIIScheduleController_1_io_valid; // @[TopModule.scala 135:15]
  assign Alu_1_io_skewing = MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_1_io_configuration = Dispatch_2_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_1_io_inputs_1 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_1_io_inputs_0 = Multiplexer_7_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_2_clock = clock;
  assign Alu_2_reset = reset;
  assign Alu_2_io_en = MultiIIScheduleController_2_io_valid; // @[TopModule.scala 135:15]
  assign Alu_2_io_skewing = MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_2_io_configuration = Dispatch_3_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_2_io_inputs_1 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_2_io_inputs_0 = Multiplexer_11_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_3_clock = clock;
  assign Alu_3_reset = reset;
  assign Alu_3_io_en = MultiIIScheduleController_3_io_valid; // @[TopModule.scala 135:15]
  assign Alu_3_io_skewing = MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_3_io_configuration = Dispatch_4_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_3_io_inputs_1 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_3_io_inputs_0 = Multiplexer_15_io_outs_0; // @[TopModule.scala 267:60]
  assign MultiIIScheduleController_clock = clock;
  assign MultiIIScheduleController_reset = reset;
  assign MultiIIScheduleController_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_io_schedules_0 = scheduleDispatch_io_outs_0; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_schedules_1 = scheduleDispatch_io_outs_1; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_schedules_2 = scheduleDispatch_io_outs_2; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_schedules_3 = scheduleDispatch_io_outs_3; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_1_clock = clock;
  assign MultiIIScheduleController_1_reset = reset;
  assign MultiIIScheduleController_1_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_1_io_schedules_0 = scheduleDispatch_io_outs_4; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_schedules_1 = scheduleDispatch_io_outs_5; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_schedules_2 = scheduleDispatch_io_outs_6; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_schedules_3 = scheduleDispatch_io_outs_7; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_2_clock = clock;
  assign MultiIIScheduleController_2_reset = reset;
  assign MultiIIScheduleController_2_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_2_io_schedules_0 = scheduleDispatch_io_outs_8; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_schedules_1 = scheduleDispatch_io_outs_9; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_schedules_2 = scheduleDispatch_io_outs_10; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_schedules_3 = scheduleDispatch_io_outs_11; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_3_clock = clock;
  assign MultiIIScheduleController_3_reset = reset;
  assign MultiIIScheduleController_3_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_3_io_schedules_0 = scheduleDispatch_io_outs_12; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_schedules_1 = scheduleDispatch_io_outs_13; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_schedules_2 = scheduleDispatch_io_outs_14; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_schedules_3 = scheduleDispatch_io_outs_15; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_II = io_II; // @[TopModule.scala 131:33]
  assign RegisterFile_clock = clock;
  assign RegisterFile_reset = reset;
  assign RegisterFile_io_configuration = Dispatch_1_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_io_inputs_0 = Alu_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_1_clock = clock;
  assign RegisterFile_1_reset = reset;
  assign RegisterFile_1_io_configuration = Dispatch_2_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_1_io_inputs_0 = Alu_1_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_2_clock = clock;
  assign RegisterFile_2_reset = reset;
  assign RegisterFile_2_io_configuration = Dispatch_3_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_2_io_inputs_0 = Alu_2_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_3_clock = clock;
  assign RegisterFile_3_reset = reset;
  assign RegisterFile_3_io_configuration = Dispatch_4_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_3_io_inputs_0 = Alu_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_io_configuration = Dispatch_io_outs_0; // @[TopModule.scala 242:22]
  assign Multiplexer_io_inputs_1 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_io_inputs_0 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_1_io_configuration = Dispatch_io_outs_1; // @[TopModule.scala 242:22]
  assign Multiplexer_1_io_inputs_1 = io_inputs_1; // @[TopModule.scala 265:60]
  assign Multiplexer_1_io_inputs_0 = io_inputs_0; // @[TopModule.scala 265:60]
  assign Multiplexer_2_io_configuration = Dispatch_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_2_io_inputs_1 = io_inputs_1; // @[TopModule.scala 265:60]
  assign Multiplexer_2_io_inputs_0 = io_inputs_0; // @[TopModule.scala 265:60]
  assign Multiplexer_3_io_configuration = Dispatch_1_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_3_io_inputs_5 = RegisterFile_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_3_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_3_io_inputs_3 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_3_io_inputs_2 = Multiplexer_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_3_io_inputs_1 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_3_io_inputs_0 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_4_io_configuration = Dispatch_1_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_4_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_4_io_inputs_3 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_4_io_inputs_2 = Multiplexer_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_4_io_inputs_1 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_4_io_inputs_0 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_configuration = Dispatch_1_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_5_io_inputs_3 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_2 = Multiplexer_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_1 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_0 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_6_io_configuration = Dispatch_1_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_6_io_inputs_1 = Multiplexer_5_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_6_io_inputs_0 = RegisterFile_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_configuration = Dispatch_2_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_7_io_inputs_5 = RegisterFile_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_4 = ConstUnit_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_3 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_2 = Multiplexer_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_1 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_0 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_8_io_configuration = Dispatch_2_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_8_io_inputs_4 = ConstUnit_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_8_io_inputs_3 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_8_io_inputs_2 = Multiplexer_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_8_io_inputs_1 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_8_io_inputs_0 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_configuration = Dispatch_2_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_9_io_inputs_3 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_2 = Multiplexer_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_1 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_0 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_10_io_configuration = Dispatch_2_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_10_io_inputs_1 = Multiplexer_9_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_10_io_inputs_0 = RegisterFile_1_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_configuration = Dispatch_3_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_11_io_inputs_5 = RegisterFile_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_4 = ConstUnit_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_3 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_2 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_1 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_0 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_12_io_configuration = Dispatch_3_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_12_io_inputs_4 = ConstUnit_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_12_io_inputs_3 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_12_io_inputs_2 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_12_io_inputs_1 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_12_io_inputs_0 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_configuration = Dispatch_3_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_13_io_inputs_3 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_2 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_1 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_0 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_14_io_configuration = Dispatch_3_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_14_io_inputs_1 = Multiplexer_13_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_14_io_inputs_0 = RegisterFile_2_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_configuration = Dispatch_4_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_15_io_inputs_5 = RegisterFile_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_4 = ConstUnit_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_3 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_2 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_1 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_0 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_16_io_configuration = Dispatch_4_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_16_io_inputs_4 = ConstUnit_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_16_io_inputs_3 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_16_io_inputs_2 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_16_io_inputs_1 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_16_io_inputs_0 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_configuration = Dispatch_4_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_17_io_inputs_3 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_2 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_1 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_0 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_18_io_configuration = Dispatch_4_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_18_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_18_io_inputs_0 = RegisterFile_3_io_outs_1; // @[TopModule.scala 267:60]
  assign ConstUnit_io_configuration = Dispatch_1_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_1_io_configuration = Dispatch_2_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_2_io_configuration = Dispatch_3_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_3_io_configuration = Dispatch_4_io_outs_6; // @[TopModule.scala 242:22]
  assign configControllers_0_clock = clock;
  assign configControllers_0_reset = reset;
  assign configControllers_0_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_0_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_0_io_inConfig = topDispatch_io_outs_0; // @[TopModule.scala 252:38]
  assign Dispatch_io_configuration = configControllers_0_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_1_clock = clock;
  assign configControllers_1_reset = reset;
  assign configControllers_1_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_1_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_1_io_inConfig = topDispatch_io_outs_1; // @[TopModule.scala 252:38]
  assign Dispatch_1_io_configuration = configControllers_1_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_2_clock = clock;
  assign configControllers_2_reset = reset;
  assign configControllers_2_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_2_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_2_io_inConfig = topDispatch_io_outs_2; // @[TopModule.scala 252:38]
  assign Dispatch_2_io_configuration = configControllers_2_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_3_clock = clock;
  assign configControllers_3_reset = reset;
  assign configControllers_3_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_3_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_3_io_inConfig = topDispatch_io_outs_3; // @[TopModule.scala 252:38]
  assign Dispatch_3_io_configuration = configControllers_3_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_4_clock = clock;
  assign configControllers_4_reset = reset;
  assign configControllers_4_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_4_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_4_io_inConfig = topDispatch_io_outs_4; // @[TopModule.scala 252:38]
  assign Dispatch_4_io_configuration = configControllers_4_io_outConfig; // @[TopModule.scala 245:31]
  assign topDispatch_io_configuration = io_configuration; // @[TopModule.scala 250:32]
endmodule
