module Dispatch(
  input  [703:0] io_configuration,
  output [10:0]  io_outs_63,
  output [10:0]  io_outs_62,
  output [10:0]  io_outs_61,
  output [10:0]  io_outs_60,
  output [10:0]  io_outs_59,
  output [10:0]  io_outs_58,
  output [10:0]  io_outs_57,
  output [10:0]  io_outs_56,
  output [10:0]  io_outs_55,
  output [10:0]  io_outs_54,
  output [10:0]  io_outs_53,
  output [10:0]  io_outs_52,
  output [10:0]  io_outs_51,
  output [10:0]  io_outs_50,
  output [10:0]  io_outs_49,
  output [10:0]  io_outs_48,
  output [10:0]  io_outs_47,
  output [10:0]  io_outs_46,
  output [10:0]  io_outs_45,
  output [10:0]  io_outs_44,
  output [10:0]  io_outs_43,
  output [10:0]  io_outs_42,
  output [10:0]  io_outs_41,
  output [10:0]  io_outs_40,
  output [10:0]  io_outs_39,
  output [10:0]  io_outs_38,
  output [10:0]  io_outs_37,
  output [10:0]  io_outs_36,
  output [10:0]  io_outs_35,
  output [10:0]  io_outs_34,
  output [10:0]  io_outs_33,
  output [10:0]  io_outs_32,
  output [10:0]  io_outs_31,
  output [10:0]  io_outs_30,
  output [10:0]  io_outs_29,
  output [10:0]  io_outs_28,
  output [10:0]  io_outs_27,
  output [10:0]  io_outs_26,
  output [10:0]  io_outs_25,
  output [10:0]  io_outs_24,
  output [10:0]  io_outs_23,
  output [10:0]  io_outs_22,
  output [10:0]  io_outs_21,
  output [10:0]  io_outs_20,
  output [10:0]  io_outs_19,
  output [10:0]  io_outs_18,
  output [10:0]  io_outs_17,
  output [10:0]  io_outs_16,
  output [10:0]  io_outs_15,
  output [10:0]  io_outs_14,
  output [10:0]  io_outs_13,
  output [10:0]  io_outs_12,
  output [10:0]  io_outs_11,
  output [10:0]  io_outs_10,
  output [10:0]  io_outs_9,
  output [10:0]  io_outs_8,
  output [10:0]  io_outs_7,
  output [10:0]  io_outs_6,
  output [10:0]  io_outs_5,
  output [10:0]  io_outs_4,
  output [10:0]  io_outs_3,
  output [10:0]  io_outs_2,
  output [10:0]  io_outs_1,
  output [10:0]  io_outs_0
);
  assign io_outs_63 = io_configuration[703:693]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_62 = io_configuration[692:682]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_61 = io_configuration[681:671]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_60 = io_configuration[670:660]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_59 = io_configuration[659:649]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_58 = io_configuration[648:638]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_57 = io_configuration[637:627]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_56 = io_configuration[626:616]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_55 = io_configuration[615:605]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_54 = io_configuration[604:594]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_53 = io_configuration[593:583]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_52 = io_configuration[582:572]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_51 = io_configuration[571:561]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_50 = io_configuration[560:550]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_49 = io_configuration[549:539]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_48 = io_configuration[538:528]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_47 = io_configuration[527:517]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_46 = io_configuration[516:506]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_45 = io_configuration[505:495]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_44 = io_configuration[494:484]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_43 = io_configuration[483:473]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_42 = io_configuration[472:462]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_41 = io_configuration[461:451]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_40 = io_configuration[450:440]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_39 = io_configuration[439:429]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_38 = io_configuration[428:418]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_37 = io_configuration[417:407]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_36 = io_configuration[406:396]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_35 = io_configuration[395:385]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_34 = io_configuration[384:374]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_33 = io_configuration[373:363]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_32 = io_configuration[362:352]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_31 = io_configuration[351:341]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_30 = io_configuration[340:330]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_29 = io_configuration[329:319]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_28 = io_configuration[318:308]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_27 = io_configuration[307:297]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_26 = io_configuration[296:286]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_25 = io_configuration[285:275]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_24 = io_configuration[274:264]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_23 = io_configuration[263:253]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_22 = io_configuration[252:242]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_21 = io_configuration[241:231]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_20 = io_configuration[230:220]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_19 = io_configuration[219:209]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_18 = io_configuration[208:198]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_17 = io_configuration[197:187]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_16 = io_configuration[186:176]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_15 = io_configuration[175:165]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_14 = io_configuration[164:154]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_13 = io_configuration[153:143]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_12 = io_configuration[142:132]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_11 = io_configuration[131:121]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_10 = io_configuration[120:110]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_9 = io_configuration[109:99]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_8 = io_configuration[98:88]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_7 = io_configuration[87:77]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_6 = io_configuration[76:66]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_5 = io_configuration[65:55]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_4 = io_configuration[54:44]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_3 = io_configuration[43:33]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_2 = io_configuration[32:22]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[21:11]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[10:0]; // @[BasicChiselModules.scala 464:18]
endmodule
module RegNextN(
  input         clock,
  input         reset,
  input  [4:0]  io_latency,
  input  [31:0] io_input,
  output [31:0] io_out
);
  reg [31:0] regArray_0; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_0;
  reg [31:0] regArray_1; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_1;
  reg [31:0] regArray_2; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_2;
  reg [31:0] regArray_3; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_3;
  reg [31:0] regArray_4; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_4;
  reg [31:0] regArray_5; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_5;
  reg [31:0] regArray_6; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_6;
  reg [31:0] regArray_7; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_7;
  reg [31:0] regArray_8; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_8;
  reg [31:0] regArray_9; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_9;
  reg [31:0] regArray_10; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_10;
  reg [31:0] regArray_11; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_11;
  reg [31:0] regArray_12; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_12;
  reg [31:0] regArray_13; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_13;
  reg [31:0] regArray_14; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_14;
  reg [31:0] regArray_15; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_15;
  reg [31:0] regArray_16; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_16;
  reg [31:0] regArray_17; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_17;
  reg [31:0] regArray_18; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_18;
  reg [31:0] regArray_19; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_19;
  reg [31:0] regArray_20; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_20;
  reg [31:0] regArray_21; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_21;
  reg [31:0] regArray_22; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_22;
  reg [31:0] regArray_23; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_23;
  reg [31:0] regArray_24; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_24;
  reg [31:0] regArray_25; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_25;
  reg [31:0] regArray_26; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_26;
  reg [31:0] regArray_27; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_27;
  reg [31:0] regArray_28; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_28;
  reg [31:0] regArray_29; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_29;
  reg [31:0] regArray_30; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_30;
  reg [31:0] regArray_31; // @[BasicChiselModules.scala 40:25]
  reg [31:0] _RAND_31;
  reg [4:0] posReg; // @[BasicChiselModules.scala 41:23]
  reg [31:0] _RAND_32;
  wire  _T_1; // @[BasicChiselModules.scala 43:19]
  wire [4:0] _T_3; // @[BasicChiselModules.scala 44:31]
  wire [31:0] _GEN_1; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_2; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_3; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_4; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_5; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_6; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_7; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_8; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_9; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_10; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_11; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_12; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_13; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_14; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_15; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_16; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_17; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_18; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_19; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_20; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_21; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_22; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_23; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_24; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_25; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_26; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_27; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_28; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_29; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_30; // @[BasicChiselModules.scala 44:12]
  wire [31:0] _GEN_31; // @[BasicChiselModules.scala 44:12]
  wire [4:0] _T_5; // @[BasicChiselModules.scala 49:20]
  assign _T_1 = io_latency > 5'h0; // @[BasicChiselModules.scala 43:19]
  assign _T_3 = posReg - io_latency; // @[BasicChiselModules.scala 44:31]
  assign _GEN_1 = 5'h1 == _T_3 ? regArray_1 : regArray_0; // @[BasicChiselModules.scala 44:12]
  assign _GEN_2 = 5'h2 == _T_3 ? regArray_2 : _GEN_1; // @[BasicChiselModules.scala 44:12]
  assign _GEN_3 = 5'h3 == _T_3 ? regArray_3 : _GEN_2; // @[BasicChiselModules.scala 44:12]
  assign _GEN_4 = 5'h4 == _T_3 ? regArray_4 : _GEN_3; // @[BasicChiselModules.scala 44:12]
  assign _GEN_5 = 5'h5 == _T_3 ? regArray_5 : _GEN_4; // @[BasicChiselModules.scala 44:12]
  assign _GEN_6 = 5'h6 == _T_3 ? regArray_6 : _GEN_5; // @[BasicChiselModules.scala 44:12]
  assign _GEN_7 = 5'h7 == _T_3 ? regArray_7 : _GEN_6; // @[BasicChiselModules.scala 44:12]
  assign _GEN_8 = 5'h8 == _T_3 ? regArray_8 : _GEN_7; // @[BasicChiselModules.scala 44:12]
  assign _GEN_9 = 5'h9 == _T_3 ? regArray_9 : _GEN_8; // @[BasicChiselModules.scala 44:12]
  assign _GEN_10 = 5'ha == _T_3 ? regArray_10 : _GEN_9; // @[BasicChiselModules.scala 44:12]
  assign _GEN_11 = 5'hb == _T_3 ? regArray_11 : _GEN_10; // @[BasicChiselModules.scala 44:12]
  assign _GEN_12 = 5'hc == _T_3 ? regArray_12 : _GEN_11; // @[BasicChiselModules.scala 44:12]
  assign _GEN_13 = 5'hd == _T_3 ? regArray_13 : _GEN_12; // @[BasicChiselModules.scala 44:12]
  assign _GEN_14 = 5'he == _T_3 ? regArray_14 : _GEN_13; // @[BasicChiselModules.scala 44:12]
  assign _GEN_15 = 5'hf == _T_3 ? regArray_15 : _GEN_14; // @[BasicChiselModules.scala 44:12]
  assign _GEN_16 = 5'h10 == _T_3 ? regArray_16 : _GEN_15; // @[BasicChiselModules.scala 44:12]
  assign _GEN_17 = 5'h11 == _T_3 ? regArray_17 : _GEN_16; // @[BasicChiselModules.scala 44:12]
  assign _GEN_18 = 5'h12 == _T_3 ? regArray_18 : _GEN_17; // @[BasicChiselModules.scala 44:12]
  assign _GEN_19 = 5'h13 == _T_3 ? regArray_19 : _GEN_18; // @[BasicChiselModules.scala 44:12]
  assign _GEN_20 = 5'h14 == _T_3 ? regArray_20 : _GEN_19; // @[BasicChiselModules.scala 44:12]
  assign _GEN_21 = 5'h15 == _T_3 ? regArray_21 : _GEN_20; // @[BasicChiselModules.scala 44:12]
  assign _GEN_22 = 5'h16 == _T_3 ? regArray_22 : _GEN_21; // @[BasicChiselModules.scala 44:12]
  assign _GEN_23 = 5'h17 == _T_3 ? regArray_23 : _GEN_22; // @[BasicChiselModules.scala 44:12]
  assign _GEN_24 = 5'h18 == _T_3 ? regArray_24 : _GEN_23; // @[BasicChiselModules.scala 44:12]
  assign _GEN_25 = 5'h19 == _T_3 ? regArray_25 : _GEN_24; // @[BasicChiselModules.scala 44:12]
  assign _GEN_26 = 5'h1a == _T_3 ? regArray_26 : _GEN_25; // @[BasicChiselModules.scala 44:12]
  assign _GEN_27 = 5'h1b == _T_3 ? regArray_27 : _GEN_26; // @[BasicChiselModules.scala 44:12]
  assign _GEN_28 = 5'h1c == _T_3 ? regArray_28 : _GEN_27; // @[BasicChiselModules.scala 44:12]
  assign _GEN_29 = 5'h1d == _T_3 ? regArray_29 : _GEN_28; // @[BasicChiselModules.scala 44:12]
  assign _GEN_30 = 5'h1e == _T_3 ? regArray_30 : _GEN_29; // @[BasicChiselModules.scala 44:12]
  assign _GEN_31 = 5'h1f == _T_3 ? regArray_31 : _GEN_30; // @[BasicChiselModules.scala 44:12]
  assign _T_5 = posReg + 5'h1; // @[BasicChiselModules.scala 49:20]
  assign io_out = _T_1 ? _GEN_31 : io_input; // @[BasicChiselModules.scala 44:12 BasicChiselModules.scala 47:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regArray_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regArray_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regArray_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regArray_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regArray_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regArray_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regArray_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regArray_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regArray_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regArray_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regArray_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regArray_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regArray_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regArray_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regArray_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regArray_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regArray_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regArray_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regArray_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regArray_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regArray_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regArray_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regArray_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regArray_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regArray_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regArray_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regArray_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regArray_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regArray_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regArray_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regArray_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regArray_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  posReg = _RAND_32[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regArray_0 <= 32'h0;
    end else if (_T_1) begin
      if (5'h0 == posReg) begin
        regArray_0 <= io_input;
      end
    end
    if (reset) begin
      regArray_1 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1 == posReg) begin
        regArray_1 <= io_input;
      end
    end
    if (reset) begin
      regArray_2 <= 32'h0;
    end else if (_T_1) begin
      if (5'h2 == posReg) begin
        regArray_2 <= io_input;
      end
    end
    if (reset) begin
      regArray_3 <= 32'h0;
    end else if (_T_1) begin
      if (5'h3 == posReg) begin
        regArray_3 <= io_input;
      end
    end
    if (reset) begin
      regArray_4 <= 32'h0;
    end else if (_T_1) begin
      if (5'h4 == posReg) begin
        regArray_4 <= io_input;
      end
    end
    if (reset) begin
      regArray_5 <= 32'h0;
    end else if (_T_1) begin
      if (5'h5 == posReg) begin
        regArray_5 <= io_input;
      end
    end
    if (reset) begin
      regArray_6 <= 32'h0;
    end else if (_T_1) begin
      if (5'h6 == posReg) begin
        regArray_6 <= io_input;
      end
    end
    if (reset) begin
      regArray_7 <= 32'h0;
    end else if (_T_1) begin
      if (5'h7 == posReg) begin
        regArray_7 <= io_input;
      end
    end
    if (reset) begin
      regArray_8 <= 32'h0;
    end else if (_T_1) begin
      if (5'h8 == posReg) begin
        regArray_8 <= io_input;
      end
    end
    if (reset) begin
      regArray_9 <= 32'h0;
    end else if (_T_1) begin
      if (5'h9 == posReg) begin
        regArray_9 <= io_input;
      end
    end
    if (reset) begin
      regArray_10 <= 32'h0;
    end else if (_T_1) begin
      if (5'ha == posReg) begin
        regArray_10 <= io_input;
      end
    end
    if (reset) begin
      regArray_11 <= 32'h0;
    end else if (_T_1) begin
      if (5'hb == posReg) begin
        regArray_11 <= io_input;
      end
    end
    if (reset) begin
      regArray_12 <= 32'h0;
    end else if (_T_1) begin
      if (5'hc == posReg) begin
        regArray_12 <= io_input;
      end
    end
    if (reset) begin
      regArray_13 <= 32'h0;
    end else if (_T_1) begin
      if (5'hd == posReg) begin
        regArray_13 <= io_input;
      end
    end
    if (reset) begin
      regArray_14 <= 32'h0;
    end else if (_T_1) begin
      if (5'he == posReg) begin
        regArray_14 <= io_input;
      end
    end
    if (reset) begin
      regArray_15 <= 32'h0;
    end else if (_T_1) begin
      if (5'hf == posReg) begin
        regArray_15 <= io_input;
      end
    end
    if (reset) begin
      regArray_16 <= 32'h0;
    end else if (_T_1) begin
      if (5'h10 == posReg) begin
        regArray_16 <= io_input;
      end
    end
    if (reset) begin
      regArray_17 <= 32'h0;
    end else if (_T_1) begin
      if (5'h11 == posReg) begin
        regArray_17 <= io_input;
      end
    end
    if (reset) begin
      regArray_18 <= 32'h0;
    end else if (_T_1) begin
      if (5'h12 == posReg) begin
        regArray_18 <= io_input;
      end
    end
    if (reset) begin
      regArray_19 <= 32'h0;
    end else if (_T_1) begin
      if (5'h13 == posReg) begin
        regArray_19 <= io_input;
      end
    end
    if (reset) begin
      regArray_20 <= 32'h0;
    end else if (_T_1) begin
      if (5'h14 == posReg) begin
        regArray_20 <= io_input;
      end
    end
    if (reset) begin
      regArray_21 <= 32'h0;
    end else if (_T_1) begin
      if (5'h15 == posReg) begin
        regArray_21 <= io_input;
      end
    end
    if (reset) begin
      regArray_22 <= 32'h0;
    end else if (_T_1) begin
      if (5'h16 == posReg) begin
        regArray_22 <= io_input;
      end
    end
    if (reset) begin
      regArray_23 <= 32'h0;
    end else if (_T_1) begin
      if (5'h17 == posReg) begin
        regArray_23 <= io_input;
      end
    end
    if (reset) begin
      regArray_24 <= 32'h0;
    end else if (_T_1) begin
      if (5'h18 == posReg) begin
        regArray_24 <= io_input;
      end
    end
    if (reset) begin
      regArray_25 <= 32'h0;
    end else if (_T_1) begin
      if (5'h19 == posReg) begin
        regArray_25 <= io_input;
      end
    end
    if (reset) begin
      regArray_26 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1a == posReg) begin
        regArray_26 <= io_input;
      end
    end
    if (reset) begin
      regArray_27 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1b == posReg) begin
        regArray_27 <= io_input;
      end
    end
    if (reset) begin
      regArray_28 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1c == posReg) begin
        regArray_28 <= io_input;
      end
    end
    if (reset) begin
      regArray_29 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1d == posReg) begin
        regArray_29 <= io_input;
      end
    end
    if (reset) begin
      regArray_30 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1e == posReg) begin
        regArray_30 <= io_input;
      end
    end
    if (reset) begin
      regArray_31 <= 32'h0;
    end else if (_T_1) begin
      if (5'h1f == posReg) begin
        regArray_31 <= io_input;
      end
    end
    if (reset) begin
      posReg <= 5'h0;
    end else begin
      posReg <= _T_5;
    end
  end
endmodule
module Synchronizer(
  input         clock,
  input         reset,
  input  [5:0]  io_skewing,
  input  [31:0] io_input0,
  input  [31:0] io_input1,
  output [31:0] io_skewedInput0,
  output [31:0] io_skewedInput1
);
  wire  regNextN_clock; // @[BasicChiselModules.scala 66:24]
  wire  regNextN_reset; // @[BasicChiselModules.scala 66:24]
  wire [4:0] regNextN_io_latency; // @[BasicChiselModules.scala 66:24]
  wire [31:0] regNextN_io_input; // @[BasicChiselModules.scala 66:24]
  wire [31:0] regNextN_io_out; // @[BasicChiselModules.scala 66:24]
  wire  signal; // @[BasicChiselModules.scala 68:26]
  RegNextN regNextN ( // @[BasicChiselModules.scala 66:24]
    .clock(regNextN_clock),
    .reset(regNextN_reset),
    .io_latency(regNextN_io_latency),
    .io_input(regNextN_io_input),
    .io_out(regNextN_io_out)
  );
  assign signal = io_skewing[5]; // @[BasicChiselModules.scala 68:26]
  assign io_skewedInput0 = signal ? regNextN_io_out : io_input0; // @[BasicChiselModules.scala 73:21 BasicChiselModules.scala 78:21]
  assign io_skewedInput1 = signal ? io_input1 : regNextN_io_out; // @[BasicChiselModules.scala 74:21 BasicChiselModules.scala 77:21]
  assign regNextN_clock = clock;
  assign regNextN_reset = reset;
  assign regNextN_io_latency = io_skewing[4:0]; // @[BasicChiselModules.scala 69:23]
  assign regNextN_io_input = signal ? io_input0 : io_input1; // @[BasicChiselModules.scala 72:23 BasicChiselModules.scala 76:23]
endmodule
module Alu(
  input         clock,
  input         reset,
  input         io_en,
  input  [5:0]  io_skewing,
  input  [3:0]  io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  synchronizer_clock; // @[BasicChiselModules.scala 242:28]
  wire  synchronizer_reset; // @[BasicChiselModules.scala 242:28]
  wire [5:0] synchronizer_io_skewing; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_input0; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_input1; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_skewedInput0; // @[BasicChiselModules.scala 242:28]
  wire [31:0] synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 242:28]
  wire [31:0] _T_1; // @[BasicChiselModules.scala 220:55]
  wire [31:0] _T_3; // @[BasicChiselModules.scala 221:55]
  wire [31:0] _T_4; // @[BasicChiselModules.scala 222:55]
  wire [31:0] _T_5; // @[BasicChiselModules.scala 223:54]
  wire [31:0] _T_6; // @[BasicChiselModules.scala 224:55]
  wire [63:0] _T_7; // @[BasicChiselModules.scala 225:55]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  wire [31:0] _T_11; // @[Mux.scala 68:16]
  wire  _T_12; // @[Mux.scala 68:19]
  wire [63:0] _T_13; // @[Mux.scala 68:16]
  wire  _T_14; // @[Mux.scala 68:19]
  wire [63:0] _T_15; // @[Mux.scala 68:16]
  wire  _T_16; // @[Mux.scala 68:19]
  wire [63:0] _T_17; // @[Mux.scala 68:16]
  wire  _T_18; // @[Mux.scala 68:19]
  wire [63:0] _T_19; // @[Mux.scala 68:16]
  wire  _T_20; // @[Mux.scala 68:19]
  wire [63:0] _T_21; // @[Mux.scala 68:16]
  wire  _T_22; // @[Mux.scala 68:19]
  wire [63:0] _T_23; // @[Mux.scala 68:16]
  wire [63:0] _GEN_0; // @[BasicChiselModules.scala 255:15]
  Synchronizer synchronizer ( // @[BasicChiselModules.scala 242:28]
    .clock(synchronizer_clock),
    .reset(synchronizer_reset),
    .io_skewing(synchronizer_io_skewing),
    .io_input0(synchronizer_io_input0),
    .io_input1(synchronizer_io_input1),
    .io_skewedInput0(synchronizer_io_skewedInput0),
    .io_skewedInput1(synchronizer_io_skewedInput1)
  );
  assign _T_1 = synchronizer_io_skewedInput0 + synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 220:55]
  assign _T_3 = synchronizer_io_skewedInput0 - synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 221:55]
  assign _T_4 = synchronizer_io_skewedInput0 & synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 222:55]
  assign _T_5 = synchronizer_io_skewedInput0 | synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 223:54]
  assign _T_6 = synchronizer_io_skewedInput0 ^ synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 224:55]
  assign _T_7 = synchronizer_io_skewedInput0 * synchronizer_io_skewedInput1; // @[BasicChiselModules.scala 225:55]
  assign _T_9 = synchronizer_io_skewedInput1; // @[Mux.scala 68:16]
  assign _T_10 = 4'hc == io_configuration; // @[Mux.scala 68:19]
  assign _T_11 = _T_10 ? synchronizer_io_skewedInput0 : _T_9; // @[Mux.scala 68:16]
  assign _T_12 = 4'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_13 = _T_12 ? _T_7 : {{32'd0}, _T_11}; // @[Mux.scala 68:16]
  assign _T_14 = 4'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_15 = _T_14 ? {{32'd0}, _T_6} : _T_13; // @[Mux.scala 68:16]
  assign _T_16 = 4'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_17 = _T_16 ? {{32'd0}, _T_5} : _T_15; // @[Mux.scala 68:16]
  assign _T_18 = 4'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_19 = _T_18 ? {{32'd0}, _T_4} : _T_17; // @[Mux.scala 68:16]
  assign _T_20 = 4'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_21 = _T_20 ? {{32'd0}, _T_3} : _T_19; // @[Mux.scala 68:16]
  assign _T_22 = 4'h0 == io_configuration; // @[Mux.scala 68:19]
  assign _T_23 = _T_22 ? {{32'd0}, _T_1} : _T_21; // @[Mux.scala 68:16]
  assign _GEN_0 = io_en ? _T_23 : 64'h0; // @[BasicChiselModules.scala 255:15]
  assign io_outs_0 = _GEN_0[31:0]; // @[BasicChiselModules.scala 256:9 BasicChiselModules.scala 259:11]
  assign synchronizer_clock = clock;
  assign synchronizer_reset = reset;
  assign synchronizer_io_skewing = io_skewing; // @[BasicChiselModules.scala 246:27]
  assign synchronizer_io_input0 = io_inputs_0; // @[BasicChiselModules.scala 243:26]
  assign synchronizer_io_input1 = io_inputs_1; // @[BasicChiselModules.scala 244:26]
endmodule
module ScheduleController(
  input        clock,
  input        reset,
  input        io_en,
  input  [4:0] io_waitCycle,
  output       io_valid
);
  reg  state; // @[BasicChiselModules.scala 139:22]
  reg [31:0] _RAND_0;
  reg [4:0] cycleReg; // @[BasicChiselModules.scala 140:21]
  reg [31:0] _RAND_1;
  wire  _T; // @[BasicChiselModules.scala 142:25]
  wire  _T_2; // @[BasicChiselModules.scala 145:16]
  wire [4:0] _T_5; // @[BasicChiselModules.scala 149:30]
  wire  _GEN_0; // @[BasicChiselModules.scala 146:39]
  wire  _GEN_2; // @[BasicChiselModules.scala 145:28]
  wire  _GEN_4; // @[BasicChiselModules.scala 144:15]
  assign _T = cycleReg == io_waitCycle; // @[BasicChiselModules.scala 142:25]
  assign _T_2 = state == 1'h0; // @[BasicChiselModules.scala 145:16]
  assign _T_5 = cycleReg + 5'h1; // @[BasicChiselModules.scala 149:30]
  assign _GEN_0 = _T | state; // @[BasicChiselModules.scala 146:39]
  assign _GEN_2 = _T_2 ? _GEN_0 : state; // @[BasicChiselModules.scala 145:28]
  assign _GEN_4 = io_en & _GEN_2; // @[BasicChiselModules.scala 144:15]
  assign io_valid = _T & io_en; // @[BasicChiselModules.scala 142:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_4;
    end
    if (io_en) begin
      if (_T_2) begin
        if (!(_T)) begin
          cycleReg <= _T_5;
        end
      end
    end else begin
      cycleReg <= 5'h0;
    end
  end
endmodule
module MultiIIScheduleController(
  input         clock,
  input         reset,
  input         io_en,
  input  [10:0] io_schedules_0,
  input  [10:0] io_schedules_1,
  input  [10:0] io_schedules_2,
  input  [10:0] io_schedules_3,
  input  [1:0]  io_II,
  output        io_valid,
  output [5:0]  io_skewing
);
  wire  ScheduleController_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_io_valid; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_1_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_1_io_valid; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_2_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_2_io_valid; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_clock; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_reset; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_io_en; // @[BasicChiselModules.scala 170:77]
  wire [4:0] ScheduleController_3_io_waitCycle; // @[BasicChiselModules.scala 170:77]
  wire  ScheduleController_3_io_valid; // @[BasicChiselModules.scala 170:77]
  reg  validRegs_0; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_0;
  reg  validRegs_1; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_1;
  reg  validRegs_2; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_2;
  reg  validRegs_3; // @[BasicChiselModules.scala 171:26]
  reg [31:0] _RAND_3;
  reg [1:0] cycleReg; // @[BasicChiselModules.scala 172:25]
  reg [31:0] _RAND_4;
  wire  _GEN_1; // @[BasicChiselModules.scala 181:12]
  wire  _GEN_2; // @[BasicChiselModules.scala 181:12]
  wire [10:0] _GEN_5; // @[BasicChiselModules.scala 182:39]
  wire [10:0] _GEN_6; // @[BasicChiselModules.scala 182:39]
  wire [10:0] _GEN_7; // @[BasicChiselModules.scala 182:39]
  wire [1:0] _T_8; // @[BasicChiselModules.scala 185:29]
  wire  _T_9; // @[BasicChiselModules.scala 185:19]
  wire [1:0] _T_11; // @[BasicChiselModules.scala 188:28]
  ScheduleController ScheduleController ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_clock),
    .reset(ScheduleController_reset),
    .io_en(ScheduleController_io_en),
    .io_waitCycle(ScheduleController_io_waitCycle),
    .io_valid(ScheduleController_io_valid)
  );
  ScheduleController ScheduleController_1 ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_1_clock),
    .reset(ScheduleController_1_reset),
    .io_en(ScheduleController_1_io_en),
    .io_waitCycle(ScheduleController_1_io_waitCycle),
    .io_valid(ScheduleController_1_io_valid)
  );
  ScheduleController ScheduleController_2 ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_2_clock),
    .reset(ScheduleController_2_reset),
    .io_en(ScheduleController_2_io_en),
    .io_waitCycle(ScheduleController_2_io_waitCycle),
    .io_valid(ScheduleController_2_io_valid)
  );
  ScheduleController ScheduleController_3 ( // @[BasicChiselModules.scala 170:77]
    .clock(ScheduleController_3_clock),
    .reset(ScheduleController_3_reset),
    .io_en(ScheduleController_3_io_en),
    .io_waitCycle(ScheduleController_3_io_waitCycle),
    .io_valid(ScheduleController_3_io_valid)
  );
  assign _GEN_1 = 2'h1 == cycleReg ? validRegs_1 : validRegs_0; // @[BasicChiselModules.scala 181:12]
  assign _GEN_2 = 2'h2 == cycleReg ? validRegs_2 : _GEN_1; // @[BasicChiselModules.scala 181:12]
  assign _GEN_5 = 2'h1 == cycleReg ? io_schedules_1 : io_schedules_0; // @[BasicChiselModules.scala 182:39]
  assign _GEN_6 = 2'h2 == cycleReg ? io_schedules_2 : _GEN_5; // @[BasicChiselModules.scala 182:39]
  assign _GEN_7 = 2'h3 == cycleReg ? io_schedules_3 : _GEN_6; // @[BasicChiselModules.scala 182:39]
  assign _T_8 = io_II - 2'h1; // @[BasicChiselModules.scala 185:29]
  assign _T_9 = cycleReg == _T_8; // @[BasicChiselModules.scala 185:19]
  assign _T_11 = cycleReg + 2'h1; // @[BasicChiselModules.scala 188:28]
  assign io_valid = 2'h3 == cycleReg ? validRegs_3 : _GEN_2; // @[BasicChiselModules.scala 181:12]
  assign io_skewing = _GEN_7[10:5]; // @[BasicChiselModules.scala 182:14]
  assign ScheduleController_clock = clock;
  assign ScheduleController_reset = reset;
  assign ScheduleController_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_io_waitCycle = io_schedules_0[4:0]; // @[BasicChiselModules.scala 177:37]
  assign ScheduleController_1_clock = clock;
  assign ScheduleController_1_reset = reset;
  assign ScheduleController_1_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_1_io_waitCycle = io_schedules_1[4:0]; // @[BasicChiselModules.scala 177:37]
  assign ScheduleController_2_clock = clock;
  assign ScheduleController_2_reset = reset;
  assign ScheduleController_2_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_2_io_waitCycle = io_schedules_2[4:0]; // @[BasicChiselModules.scala 177:37]
  assign ScheduleController_3_clock = clock;
  assign ScheduleController_3_reset = reset;
  assign ScheduleController_3_io_en = io_en; // @[BasicChiselModules.scala 176:30]
  assign ScheduleController_3_io_waitCycle = io_schedules_3[4:0]; // @[BasicChiselModules.scala 177:37]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validRegs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  validRegs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  validRegs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  validRegs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cycleReg = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      validRegs_0 <= 1'h0;
    end else begin
      validRegs_0 <= ScheduleController_io_valid;
    end
    if (reset) begin
      validRegs_1 <= 1'h0;
    end else begin
      validRegs_1 <= ScheduleController_1_io_valid;
    end
    if (reset) begin
      validRegs_2 <= 1'h0;
    end else begin
      validRegs_2 <= ScheduleController_2_io_valid;
    end
    if (reset) begin
      validRegs_3 <= 1'h0;
    end else begin
      validRegs_3 <= ScheduleController_3_io_valid;
    end
    if (reset) begin
      cycleReg <= 2'h3;
    end else if (io_en) begin
      if (_T_9) begin
        cycleReg <= 2'h0;
      end else begin
        cycleReg <= _T_11;
      end
    end
  end
endmodule
module Dispatch_1(
  input  [2:0] io_configuration,
  output       io_outs_2,
  output       io_outs_1,
  output       io_outs_0
);
  assign io_outs_2 = io_configuration[2]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[1]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[0]; // @[BasicChiselModules.scala 464:18]
endmodule
module RegisterFile(
  input         clock,
  input         reset,
  input  [3:0]  io_configuration,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_1,
  output [31:0] io_outs_0
);
  wire [2:0] Dispatch_io_configuration; // @[BasicChiselModules.scala 332:26]
  wire  Dispatch_io_outs_2; // @[BasicChiselModules.scala 332:26]
  wire  Dispatch_io_outs_1; // @[BasicChiselModules.scala 332:26]
  wire  Dispatch_io_outs_0; // @[BasicChiselModules.scala 332:26]
  wire  _T_1; // @[BasicChiselModules.scala 336:37]
  reg [31:0] _T_3_0; // @[BasicChiselModules.scala 338:23]
  reg [31:0] _RAND_0;
  reg [31:0] _T_3_1; // @[BasicChiselModules.scala 338:23]
  reg [31:0] _RAND_1;
  wire  _T_4; // @[BasicChiselModules.scala 340:20]
  Dispatch_1 Dispatch ( // @[BasicChiselModules.scala 332:26]
    .io_configuration(Dispatch_io_configuration),
    .io_outs_2(Dispatch_io_outs_2),
    .io_outs_1(Dispatch_io_outs_1),
    .io_outs_0(Dispatch_io_outs_0)
  );
  assign _T_1 = io_configuration[3]; // @[BasicChiselModules.scala 336:37]
  assign _T_4 = _T_1 == 1'h0; // @[BasicChiselModules.scala 340:20]
  assign io_outs_1 = Dispatch_io_outs_2 ? _T_3_1 : _T_3_0; // @[BasicChiselModules.scala 346:18]
  assign io_outs_0 = Dispatch_io_outs_1 ? _T_3_1 : _T_3_0; // @[BasicChiselModules.scala 346:18]
  assign Dispatch_io_configuration = io_configuration[2:0]; // @[BasicChiselModules.scala 334:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3_0 <= 32'h0;
    end else if (_T_4) begin
      if (1'h0 == Dispatch_io_outs_0) begin
        _T_3_0 <= io_inputs_0;
      end
    end
    if (reset) begin
      _T_3_1 <= 32'h0;
    end else if (_T_4) begin
      if (Dispatch_io_outs_0) begin
        _T_3_1 <= io_inputs_0;
      end
    end
  end
endmodule
module Multiplexer(
  input  [1:0]  io_configuration,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  assign _T = 2'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_3 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 2'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_2 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 2'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_1 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 2'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_6 ? io_inputs_0 : _T_5; // @[BasicChiselModules.scala 370:14]
endmodule
module Multiplexer_1(
  input         io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  assign _T_1 = io_configuration ? io_inputs_1 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 1'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_2 ? io_inputs_0 : _T_1; // @[BasicChiselModules.scala 370:14]
endmodule
module Multiplexer_5(
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_5,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  assign _T = 3'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_5 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_4 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_3 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_2 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_9 = _T_8 ? io_inputs_1 : _T_7; // @[Mux.scala 68:16]
  assign _T_10 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_10 ? io_inputs_0 : _T_9; // @[BasicChiselModules.scala 370:14]
endmodule
module Multiplexer_6(
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  assign _T = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_4 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_3 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_2 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_1 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign io_outs_0 = _T_8 ? io_inputs_0 : _T_7; // @[BasicChiselModules.scala 370:14]
endmodule
module ConstUnit(
  input  [31:0] io_configuration,
  output [31:0] io_outs_0
);
  assign io_outs_0 = io_configuration; // @[BasicChiselModules.scala 403:14]
endmodule
module ConfigController(
  input        clock,
  input        reset,
  input        io_en,
  input  [1:0] io_II,
  input  [5:0] io_inConfig,
  output [5:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 96:22]
  reg [31:0] _RAND_0;
  reg [1:0] cycleReg; // @[BasicChiselModules.scala 97:21]
  reg [31:0] _RAND_1;
  reg [5:0] configRegs_0; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_2;
  reg [5:0] configRegs_1; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_3;
  reg [5:0] configRegs_2; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_4;
  reg [5:0] configRegs_3; // @[BasicChiselModules.scala 99:27]
  reg [31:0] _RAND_5;
  wire  _T_1; // @[BasicChiselModules.scala 103:14]
  wire [5:0] _GEN_1; // @[BasicChiselModules.scala 106:18]
  wire [5:0] _GEN_2; // @[BasicChiselModules.scala 106:18]
  wire [5:0] _GEN_3; // @[BasicChiselModules.scala 106:18]
  wire  _T_3; // @[BasicChiselModules.scala 112:21]
  wire [1:0] _T_5; // @[BasicChiselModules.scala 116:30]
  wire  _GEN_9; // @[BasicChiselModules.scala 112:32]
  wire [1:0] _T_7; // @[BasicChiselModules.scala 119:31]
  wire  _T_8; // @[BasicChiselModules.scala 119:21]
  wire  _GEN_16; // @[BasicChiselModules.scala 110:34]
  wire  _GEN_22; // @[BasicChiselModules.scala 109:15]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 103:14]
  assign _GEN_1 = 2'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 106:18]
  assign _GEN_2 = 2'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 106:18]
  assign _GEN_3 = 2'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 106:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 112:21]
  assign _T_5 = cycleReg + 2'h1; // @[BasicChiselModules.scala 116:30]
  assign _GEN_9 = _T_3 | state; // @[BasicChiselModules.scala 112:32]
  assign _T_7 = io_II - 2'h1; // @[BasicChiselModules.scala 119:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 119:21]
  assign _GEN_16 = _T_1 ? _GEN_9 : state; // @[BasicChiselModules.scala 110:34]
  assign _GEN_22 = io_en & _GEN_16; // @[BasicChiselModules.scala 109:15]
  assign io_outConfig = _T_1 ? 6'h0 : _GEN_3; // @[BasicChiselModules.scala 104:18 BasicChiselModules.scala 106:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  configRegs_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  configRegs_1 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  configRegs_2 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  configRegs_3 = _RAND_5[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_22;
    end
    if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 2'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 2'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 2'h0;
    end
    if (reset) begin
      configRegs_0 <= 6'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h0 == cycleReg) begin
          configRegs_0 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 6'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h1 == cycleReg) begin
          configRegs_1 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 6'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h2 == cycleReg) begin
          configRegs_2 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 6'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h3 == cycleReg) begin
          configRegs_3 <= io_inConfig;
        end
      end
    end
  end
endmodule
module Dispatch_17(
  input  [5:0] io_configuration,
  output       io_outs_4,
  output       io_outs_3,
  output       io_outs_2,
  output       io_outs_1,
  output [1:0] io_outs_0
);
  assign io_outs_4 = io_configuration[5]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_3 = io_configuration[4]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_2 = io_configuration[3]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[2]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[1:0]; // @[BasicChiselModules.scala 464:18]
endmodule
module ConfigController_1(
  input         clock,
  input         reset,
  input         io_en,
  input  [1:0]  io_II,
  input  [48:0] io_inConfig,
  output [48:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 96:22]
  reg [31:0] _RAND_0;
  reg [1:0] cycleReg; // @[BasicChiselModules.scala 97:21]
  reg [31:0] _RAND_1;
  reg [48:0] configRegs_0; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_2;
  reg [48:0] configRegs_1; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_3;
  reg [48:0] configRegs_2; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_4;
  reg [48:0] configRegs_3; // @[BasicChiselModules.scala 99:27]
  reg [63:0] _RAND_5;
  wire  _T_1; // @[BasicChiselModules.scala 103:14]
  wire [48:0] _GEN_1; // @[BasicChiselModules.scala 106:18]
  wire [48:0] _GEN_2; // @[BasicChiselModules.scala 106:18]
  wire [48:0] _GEN_3; // @[BasicChiselModules.scala 106:18]
  wire  _T_3; // @[BasicChiselModules.scala 112:21]
  wire [1:0] _T_5; // @[BasicChiselModules.scala 116:30]
  wire  _GEN_9; // @[BasicChiselModules.scala 112:32]
  wire [1:0] _T_7; // @[BasicChiselModules.scala 119:31]
  wire  _T_8; // @[BasicChiselModules.scala 119:21]
  wire  _GEN_16; // @[BasicChiselModules.scala 110:34]
  wire  _GEN_22; // @[BasicChiselModules.scala 109:15]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 103:14]
  assign _GEN_1 = 2'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 106:18]
  assign _GEN_2 = 2'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 106:18]
  assign _GEN_3 = 2'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 106:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 112:21]
  assign _T_5 = cycleReg + 2'h1; // @[BasicChiselModules.scala 116:30]
  assign _GEN_9 = _T_3 | state; // @[BasicChiselModules.scala 112:32]
  assign _T_7 = io_II - 2'h1; // @[BasicChiselModules.scala 119:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 119:21]
  assign _GEN_16 = _T_1 ? _GEN_9 : state; // @[BasicChiselModules.scala 110:34]
  assign _GEN_22 = io_en & _GEN_16; // @[BasicChiselModules.scala 109:15]
  assign io_outConfig = _T_1 ? 49'h0 : _GEN_3; // @[BasicChiselModules.scala 104:18 BasicChiselModules.scala 106:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  configRegs_0 = _RAND_2[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  configRegs_1 = _RAND_3[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  configRegs_2 = _RAND_4[48:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  configRegs_3 = _RAND_5[48:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_22;
    end
    if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 2'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 2'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 2'h0;
    end
    if (reset) begin
      configRegs_0 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h0 == cycleReg) begin
          configRegs_0 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h1 == cycleReg) begin
          configRegs_1 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h2 == cycleReg) begin
          configRegs_2 <= io_inConfig;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 49'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (2'h3 == cycleReg) begin
          configRegs_3 <= io_inConfig;
        end
      end
    end
  end
endmodule
module Dispatch_18(
  input  [48:0] io_configuration,
  output [31:0] io_outs_6,
  output        io_outs_5,
  output [1:0]  io_outs_4,
  output [2:0]  io_outs_3,
  output [2:0]  io_outs_2,
  output [3:0]  io_outs_1,
  output [3:0]  io_outs_0
);
  assign io_outs_6 = io_configuration[48:17]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_5 = io_configuration[16]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_4 = io_configuration[15:14]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_3 = io_configuration[13:11]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_2 = io_configuration[10:8]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[7:4]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[3:0]; // @[BasicChiselModules.scala 464:18]
endmodule
module Dispatch_34(
  input  [789:0] io_configuration,
  output [48:0]  io_outs_16,
  output [48:0]  io_outs_15,
  output [48:0]  io_outs_14,
  output [48:0]  io_outs_13,
  output [48:0]  io_outs_12,
  output [48:0]  io_outs_11,
  output [48:0]  io_outs_10,
  output [48:0]  io_outs_9,
  output [48:0]  io_outs_8,
  output [48:0]  io_outs_7,
  output [48:0]  io_outs_6,
  output [48:0]  io_outs_5,
  output [48:0]  io_outs_4,
  output [48:0]  io_outs_3,
  output [48:0]  io_outs_2,
  output [48:0]  io_outs_1,
  output [5:0]   io_outs_0
);
  assign io_outs_16 = io_configuration[789:741]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_15 = io_configuration[740:692]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_14 = io_configuration[691:643]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_13 = io_configuration[642:594]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_12 = io_configuration[593:545]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_11 = io_configuration[544:496]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_10 = io_configuration[495:447]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_9 = io_configuration[446:398]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_8 = io_configuration[397:349]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_7 = io_configuration[348:300]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_6 = io_configuration[299:251]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_5 = io_configuration[250:202]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_4 = io_configuration[201:153]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_3 = io_configuration[152:104]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_2 = io_configuration[103:55]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_1 = io_configuration[54:6]; // @[BasicChiselModules.scala 464:18]
  assign io_outs_0 = io_configuration[5:0]; // @[BasicChiselModules.scala 464:18]
endmodule
module TopModule(
  input          clock,
  input          reset,
  input          io_enConfig,
  input          io_en,
  input  [703:0] io_schedules,
  input  [1:0]   io_II,
  input  [789:0] io_configuration,
  input  [31:0]  io_inputs_1,
  input  [31:0]  io_inputs_0,
  output [31:0]  io_outs_0
);
  wire [703:0] scheduleDispatch_io_configuration; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_63; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_62; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_61; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_60; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_59; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_58; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_57; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_56; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_55; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_54; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_53; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_52; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_51; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_50; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_49; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_48; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_47; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_46; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_45; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_44; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_43; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_42; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_41; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_40; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_39; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_38; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_37; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_36; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_35; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_34; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_33; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_32; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_31; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_30; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_29; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_28; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_27; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_26; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_25; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_24; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_23; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_22; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_21; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_20; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_19; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_18; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_17; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_16; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_15; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_14; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_13; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_12; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_11; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_10; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_9; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_8; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_7; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_6; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_5; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_4; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_3; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_2; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_1; // @[TopModule.scala 119:32]
  wire [10:0] scheduleDispatch_io_outs_0; // @[TopModule.scala 119:32]
  wire  Alu_clock; // @[TopModule.scala 124:54]
  wire  Alu_reset; // @[TopModule.scala 124:54]
  wire  Alu_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_1_clock; // @[TopModule.scala 124:54]
  wire  Alu_1_reset; // @[TopModule.scala 124:54]
  wire  Alu_1_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_1_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_1_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_1_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_1_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_1_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_2_clock; // @[TopModule.scala 124:54]
  wire  Alu_2_reset; // @[TopModule.scala 124:54]
  wire  Alu_2_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_2_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_2_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_2_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_2_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_2_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_3_clock; // @[TopModule.scala 124:54]
  wire  Alu_3_reset; // @[TopModule.scala 124:54]
  wire  Alu_3_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_3_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_3_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_3_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_3_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_3_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_4_clock; // @[TopModule.scala 124:54]
  wire  Alu_4_reset; // @[TopModule.scala 124:54]
  wire  Alu_4_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_4_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_4_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_4_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_4_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_4_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_5_clock; // @[TopModule.scala 124:54]
  wire  Alu_5_reset; // @[TopModule.scala 124:54]
  wire  Alu_5_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_5_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_5_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_5_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_5_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_5_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_6_clock; // @[TopModule.scala 124:54]
  wire  Alu_6_reset; // @[TopModule.scala 124:54]
  wire  Alu_6_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_6_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_6_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_6_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_6_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_6_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_7_clock; // @[TopModule.scala 124:54]
  wire  Alu_7_reset; // @[TopModule.scala 124:54]
  wire  Alu_7_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_7_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_7_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_7_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_7_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_7_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_8_clock; // @[TopModule.scala 124:54]
  wire  Alu_8_reset; // @[TopModule.scala 124:54]
  wire  Alu_8_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_8_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_8_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_8_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_8_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_8_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_9_clock; // @[TopModule.scala 124:54]
  wire  Alu_9_reset; // @[TopModule.scala 124:54]
  wire  Alu_9_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_9_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_9_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_9_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_9_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_9_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_10_clock; // @[TopModule.scala 124:54]
  wire  Alu_10_reset; // @[TopModule.scala 124:54]
  wire  Alu_10_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_10_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_10_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_10_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_10_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_10_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_11_clock; // @[TopModule.scala 124:54]
  wire  Alu_11_reset; // @[TopModule.scala 124:54]
  wire  Alu_11_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_11_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_11_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_11_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_11_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_11_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_12_clock; // @[TopModule.scala 124:54]
  wire  Alu_12_reset; // @[TopModule.scala 124:54]
  wire  Alu_12_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_12_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_12_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_12_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_12_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_12_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_13_clock; // @[TopModule.scala 124:54]
  wire  Alu_13_reset; // @[TopModule.scala 124:54]
  wire  Alu_13_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_13_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_13_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_13_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_13_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_13_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_14_clock; // @[TopModule.scala 124:54]
  wire  Alu_14_reset; // @[TopModule.scala 124:54]
  wire  Alu_14_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_14_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_14_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_14_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_14_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_14_io_outs_0; // @[TopModule.scala 124:54]
  wire  Alu_15_clock; // @[TopModule.scala 124:54]
  wire  Alu_15_reset; // @[TopModule.scala 124:54]
  wire  Alu_15_io_en; // @[TopModule.scala 124:54]
  wire [5:0] Alu_15_io_skewing; // @[TopModule.scala 124:54]
  wire [3:0] Alu_15_io_configuration; // @[TopModule.scala 124:54]
  wire [31:0] Alu_15_io_inputs_1; // @[TopModule.scala 124:54]
  wire [31:0] Alu_15_io_inputs_0; // @[TopModule.scala 124:54]
  wire [31:0] Alu_15_io_outs_0; // @[TopModule.scala 124:54]
  wire  MultiIIScheduleController_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_1_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_1_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_1_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_2_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_2_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_2_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_3_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_3_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_3_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_4_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_4_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_4_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_4_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_4_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_4_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_4_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_4_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_4_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_4_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_5_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_5_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_5_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_5_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_5_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_5_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_5_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_5_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_5_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_5_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_6_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_6_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_6_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_6_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_6_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_6_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_6_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_6_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_6_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_6_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_7_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_7_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_7_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_7_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_7_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_7_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_7_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_7_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_7_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_7_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_8_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_8_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_8_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_8_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_8_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_8_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_8_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_8_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_8_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_8_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_9_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_9_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_9_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_9_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_9_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_9_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_9_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_9_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_9_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_9_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_10_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_10_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_10_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_10_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_10_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_10_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_10_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_10_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_10_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_10_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_11_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_11_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_11_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_11_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_11_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_11_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_11_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_11_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_11_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_11_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_12_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_12_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_12_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_12_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_12_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_12_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_12_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_12_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_12_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_12_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_13_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_13_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_13_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_13_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_13_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_13_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_13_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_13_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_13_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_13_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_14_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_14_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_14_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_14_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_14_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_14_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_14_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_14_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_14_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_14_io_skewing; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_15_clock; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_15_reset; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_15_io_en; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_15_io_schedules_0; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_15_io_schedules_1; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_15_io_schedules_2; // @[TopModule.scala 126:72]
  wire [10:0] MultiIIScheduleController_15_io_schedules_3; // @[TopModule.scala 126:72]
  wire [1:0] MultiIIScheduleController_15_io_II; // @[TopModule.scala 126:72]
  wire  MultiIIScheduleController_15_io_valid; // @[TopModule.scala 126:72]
  wire [5:0] MultiIIScheduleController_15_io_skewing; // @[TopModule.scala 126:72]
  wire  RegisterFile_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_1_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_1_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_1_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_1_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_1_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_1_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_2_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_2_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_2_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_2_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_2_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_2_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_3_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_3_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_3_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_3_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_3_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_3_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_4_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_4_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_4_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_4_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_4_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_4_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_5_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_5_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_5_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_5_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_5_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_5_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_6_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_6_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_6_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_6_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_6_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_6_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_7_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_7_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_7_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_7_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_7_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_7_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_8_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_8_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_8_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_8_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_8_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_8_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_9_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_9_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_9_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_9_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_9_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_9_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_10_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_10_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_10_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_10_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_10_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_10_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_11_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_11_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_11_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_11_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_11_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_11_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_12_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_12_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_12_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_12_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_12_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_12_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_13_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_13_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_13_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_13_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_13_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_13_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_14_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_14_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_14_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_14_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_14_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_14_io_outs_0; // @[TopModule.scala 142:21]
  wire  RegisterFile_15_clock; // @[TopModule.scala 142:21]
  wire  RegisterFile_15_reset; // @[TopModule.scala 142:21]
  wire [3:0] RegisterFile_15_io_configuration; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_15_io_inputs_0; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_15_io_outs_1; // @[TopModule.scala 142:21]
  wire [31:0] RegisterFile_15_io_outs_0; // @[TopModule.scala 142:21]
  wire [1:0] Multiplexer_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_1_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_1_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_1_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_1_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_2_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_2_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_2_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_2_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_3_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_3_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_4_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_4_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_5_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_5_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_6_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_6_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_7_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_7_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_8_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_8_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_9_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_9_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_10_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_10_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_11_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_11_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_12_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_12_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_13_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_13_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_14_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_14_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_15_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_15_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_16_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_16_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_17_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_17_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_18_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_18_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_19_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_19_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_19_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_19_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_19_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_19_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_20_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_20_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_20_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_20_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_21_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_21_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_21_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_21_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_21_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_21_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_21_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_21_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_22_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_22_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_22_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_22_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_22_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_22_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_22_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_23_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_23_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_23_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_23_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_23_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_23_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_24_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_24_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_24_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_24_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_25_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_25_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_25_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_25_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_25_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_25_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_25_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_25_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_26_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_26_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_26_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_26_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_26_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_26_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_26_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_27_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_27_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_27_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_27_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_27_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_27_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_28_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_28_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_28_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_28_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_29_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_29_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_29_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_29_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_29_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_29_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_29_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_29_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_30_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_30_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_30_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_30_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_30_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_30_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_30_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_31_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_31_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_31_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_31_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_31_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_31_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_32_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_32_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_32_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_32_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_33_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_33_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_33_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_33_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_33_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_33_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_33_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_33_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_34_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_34_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_34_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_34_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_34_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_34_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_34_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_35_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_35_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_35_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_35_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_35_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_35_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_36_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_36_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_36_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_36_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_37_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_37_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_37_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_37_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_37_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_37_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_37_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_37_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_38_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_38_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_38_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_38_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_38_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_38_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_38_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_39_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_39_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_39_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_39_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_39_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_39_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_40_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_40_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_40_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_40_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_41_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_41_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_41_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_41_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_41_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_41_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_41_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_41_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_42_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_42_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_42_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_42_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_42_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_42_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_42_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_43_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_43_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_43_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_43_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_43_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_43_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_44_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_44_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_44_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_44_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_45_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_45_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_45_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_45_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_45_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_45_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_45_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_45_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_46_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_46_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_46_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_46_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_46_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_46_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_46_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_47_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_47_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_47_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_47_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_47_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_47_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_48_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_48_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_48_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_48_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_49_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_49_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_49_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_49_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_49_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_49_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_49_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_49_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_50_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_50_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_50_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_50_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_50_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_50_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_50_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_51_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_51_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_51_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_51_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_51_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_51_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_52_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_52_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_52_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_52_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_53_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_53_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_53_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_53_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_53_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_53_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_53_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_53_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_54_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_54_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_54_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_54_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_54_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_54_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_54_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_55_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_55_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_55_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_55_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_55_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_55_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_56_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_56_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_56_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_56_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_57_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_57_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_57_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_57_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_57_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_57_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_57_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_57_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_58_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_58_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_58_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_58_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_58_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_58_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_58_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_59_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_59_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_59_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_59_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_59_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_59_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_60_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_60_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_60_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_60_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_61_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_61_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_61_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_61_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_61_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_61_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_61_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_61_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_62_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_62_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_62_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_62_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_62_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_62_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_62_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_63_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_63_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_63_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_63_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_63_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_63_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_64_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_64_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_64_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_64_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_65_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_65_io_inputs_5; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_65_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_65_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_65_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_65_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_65_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_65_io_outs_0; // @[TopModule.scala 153:11]
  wire [2:0] Multiplexer_66_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_66_io_inputs_4; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_66_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_66_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_66_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_66_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_66_io_outs_0; // @[TopModule.scala 153:11]
  wire [1:0] Multiplexer_67_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_67_io_inputs_3; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_67_io_inputs_2; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_67_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_67_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_67_io_outs_0; // @[TopModule.scala 153:11]
  wire  Multiplexer_68_io_configuration; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_68_io_inputs_1; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_68_io_inputs_0; // @[TopModule.scala 153:11]
  wire [31:0] Multiplexer_68_io_outs_0; // @[TopModule.scala 153:11]
  wire [31:0] ConstUnit_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_1_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_1_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_2_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_2_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_3_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_3_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_4_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_4_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_5_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_5_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_6_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_6_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_7_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_7_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_8_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_8_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_9_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_9_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_10_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_10_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_11_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_11_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_12_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_12_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_13_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_13_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_14_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_14_io_outs_0; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_15_io_configuration; // @[TopModule.scala 161:21]
  wire [31:0] ConstUnit_15_io_outs_0; // @[TopModule.scala 161:21]
  wire  configControllers_0_clock; // @[TopModule.scala 234:34]
  wire  configControllers_0_reset; // @[TopModule.scala 234:34]
  wire  configControllers_0_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_0_io_II; // @[TopModule.scala 234:34]
  wire [5:0] configControllers_0_io_inConfig; // @[TopModule.scala 234:34]
  wire [5:0] configControllers_0_io_outConfig; // @[TopModule.scala 234:34]
  wire [5:0] Dispatch_io_configuration; // @[TopModule.scala 239:26]
  wire  Dispatch_io_outs_4; // @[TopModule.scala 239:26]
  wire  Dispatch_io_outs_3; // @[TopModule.scala 239:26]
  wire  Dispatch_io_outs_2; // @[TopModule.scala 239:26]
  wire  Dispatch_io_outs_1; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_1_clock; // @[TopModule.scala 234:34]
  wire  configControllers_1_reset; // @[TopModule.scala 234:34]
  wire  configControllers_1_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_1_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_1_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_1_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_1_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_1_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_1_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_1_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_1_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_1_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_1_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_1_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_2_clock; // @[TopModule.scala 234:34]
  wire  configControllers_2_reset; // @[TopModule.scala 234:34]
  wire  configControllers_2_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_2_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_2_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_2_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_2_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_2_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_2_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_2_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_2_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_2_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_2_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_2_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_3_clock; // @[TopModule.scala 234:34]
  wire  configControllers_3_reset; // @[TopModule.scala 234:34]
  wire  configControllers_3_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_3_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_3_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_3_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_3_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_3_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_3_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_3_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_3_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_3_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_3_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_3_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_4_clock; // @[TopModule.scala 234:34]
  wire  configControllers_4_reset; // @[TopModule.scala 234:34]
  wire  configControllers_4_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_4_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_4_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_4_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_4_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_4_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_4_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_4_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_4_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_4_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_4_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_4_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_5_clock; // @[TopModule.scala 234:34]
  wire  configControllers_5_reset; // @[TopModule.scala 234:34]
  wire  configControllers_5_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_5_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_5_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_5_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_5_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_5_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_5_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_5_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_5_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_5_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_5_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_5_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_6_clock; // @[TopModule.scala 234:34]
  wire  configControllers_6_reset; // @[TopModule.scala 234:34]
  wire  configControllers_6_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_6_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_6_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_6_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_6_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_6_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_6_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_6_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_6_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_6_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_6_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_6_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_7_clock; // @[TopModule.scala 234:34]
  wire  configControllers_7_reset; // @[TopModule.scala 234:34]
  wire  configControllers_7_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_7_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_7_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_7_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_7_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_7_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_7_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_7_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_7_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_7_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_7_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_7_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_8_clock; // @[TopModule.scala 234:34]
  wire  configControllers_8_reset; // @[TopModule.scala 234:34]
  wire  configControllers_8_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_8_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_8_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_8_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_8_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_8_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_8_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_8_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_8_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_8_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_8_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_8_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_9_clock; // @[TopModule.scala 234:34]
  wire  configControllers_9_reset; // @[TopModule.scala 234:34]
  wire  configControllers_9_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_9_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_9_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_9_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_9_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_9_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_9_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_9_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_9_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_9_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_9_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_9_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_10_clock; // @[TopModule.scala 234:34]
  wire  configControllers_10_reset; // @[TopModule.scala 234:34]
  wire  configControllers_10_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_10_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_10_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_10_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_10_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_10_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_10_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_10_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_10_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_10_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_10_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_10_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_11_clock; // @[TopModule.scala 234:34]
  wire  configControllers_11_reset; // @[TopModule.scala 234:34]
  wire  configControllers_11_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_11_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_11_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_11_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_11_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_11_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_11_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_11_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_11_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_11_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_11_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_11_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_12_clock; // @[TopModule.scala 234:34]
  wire  configControllers_12_reset; // @[TopModule.scala 234:34]
  wire  configControllers_12_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_12_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_12_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_12_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_12_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_12_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_12_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_12_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_12_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_12_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_12_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_12_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_13_clock; // @[TopModule.scala 234:34]
  wire  configControllers_13_reset; // @[TopModule.scala 234:34]
  wire  configControllers_13_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_13_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_13_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_13_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_13_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_13_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_13_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_13_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_13_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_13_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_13_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_13_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_14_clock; // @[TopModule.scala 234:34]
  wire  configControllers_14_reset; // @[TopModule.scala 234:34]
  wire  configControllers_14_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_14_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_14_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_14_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_14_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_14_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_14_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_14_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_14_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_14_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_14_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_14_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_15_clock; // @[TopModule.scala 234:34]
  wire  configControllers_15_reset; // @[TopModule.scala 234:34]
  wire  configControllers_15_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_15_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_15_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_15_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_15_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_15_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_15_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_15_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_15_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_15_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_15_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_15_io_outs_0; // @[TopModule.scala 239:26]
  wire  configControllers_16_clock; // @[TopModule.scala 234:34]
  wire  configControllers_16_reset; // @[TopModule.scala 234:34]
  wire  configControllers_16_io_en; // @[TopModule.scala 234:34]
  wire [1:0] configControllers_16_io_II; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_16_io_inConfig; // @[TopModule.scala 234:34]
  wire [48:0] configControllers_16_io_outConfig; // @[TopModule.scala 234:34]
  wire [48:0] Dispatch_16_io_configuration; // @[TopModule.scala 239:26]
  wire [31:0] Dispatch_16_io_outs_6; // @[TopModule.scala 239:26]
  wire  Dispatch_16_io_outs_5; // @[TopModule.scala 239:26]
  wire [1:0] Dispatch_16_io_outs_4; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_16_io_outs_3; // @[TopModule.scala 239:26]
  wire [2:0] Dispatch_16_io_outs_2; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_16_io_outs_1; // @[TopModule.scala 239:26]
  wire [3:0] Dispatch_16_io_outs_0; // @[TopModule.scala 239:26]
  wire [789:0] topDispatch_io_configuration; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_16; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_15; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_14; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_13; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_12; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_11; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_10; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_9; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_8; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_7; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_6; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_5; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_4; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_3; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_2; // @[TopModule.scala 248:27]
  wire [48:0] topDispatch_io_outs_1; // @[TopModule.scala 248:27]
  wire [5:0] topDispatch_io_outs_0; // @[TopModule.scala 248:27]
  Dispatch scheduleDispatch ( // @[TopModule.scala 119:32]
    .io_configuration(scheduleDispatch_io_configuration),
    .io_outs_63(scheduleDispatch_io_outs_63),
    .io_outs_62(scheduleDispatch_io_outs_62),
    .io_outs_61(scheduleDispatch_io_outs_61),
    .io_outs_60(scheduleDispatch_io_outs_60),
    .io_outs_59(scheduleDispatch_io_outs_59),
    .io_outs_58(scheduleDispatch_io_outs_58),
    .io_outs_57(scheduleDispatch_io_outs_57),
    .io_outs_56(scheduleDispatch_io_outs_56),
    .io_outs_55(scheduleDispatch_io_outs_55),
    .io_outs_54(scheduleDispatch_io_outs_54),
    .io_outs_53(scheduleDispatch_io_outs_53),
    .io_outs_52(scheduleDispatch_io_outs_52),
    .io_outs_51(scheduleDispatch_io_outs_51),
    .io_outs_50(scheduleDispatch_io_outs_50),
    .io_outs_49(scheduleDispatch_io_outs_49),
    .io_outs_48(scheduleDispatch_io_outs_48),
    .io_outs_47(scheduleDispatch_io_outs_47),
    .io_outs_46(scheduleDispatch_io_outs_46),
    .io_outs_45(scheduleDispatch_io_outs_45),
    .io_outs_44(scheduleDispatch_io_outs_44),
    .io_outs_43(scheduleDispatch_io_outs_43),
    .io_outs_42(scheduleDispatch_io_outs_42),
    .io_outs_41(scheduleDispatch_io_outs_41),
    .io_outs_40(scheduleDispatch_io_outs_40),
    .io_outs_39(scheduleDispatch_io_outs_39),
    .io_outs_38(scheduleDispatch_io_outs_38),
    .io_outs_37(scheduleDispatch_io_outs_37),
    .io_outs_36(scheduleDispatch_io_outs_36),
    .io_outs_35(scheduleDispatch_io_outs_35),
    .io_outs_34(scheduleDispatch_io_outs_34),
    .io_outs_33(scheduleDispatch_io_outs_33),
    .io_outs_32(scheduleDispatch_io_outs_32),
    .io_outs_31(scheduleDispatch_io_outs_31),
    .io_outs_30(scheduleDispatch_io_outs_30),
    .io_outs_29(scheduleDispatch_io_outs_29),
    .io_outs_28(scheduleDispatch_io_outs_28),
    .io_outs_27(scheduleDispatch_io_outs_27),
    .io_outs_26(scheduleDispatch_io_outs_26),
    .io_outs_25(scheduleDispatch_io_outs_25),
    .io_outs_24(scheduleDispatch_io_outs_24),
    .io_outs_23(scheduleDispatch_io_outs_23),
    .io_outs_22(scheduleDispatch_io_outs_22),
    .io_outs_21(scheduleDispatch_io_outs_21),
    .io_outs_20(scheduleDispatch_io_outs_20),
    .io_outs_19(scheduleDispatch_io_outs_19),
    .io_outs_18(scheduleDispatch_io_outs_18),
    .io_outs_17(scheduleDispatch_io_outs_17),
    .io_outs_16(scheduleDispatch_io_outs_16),
    .io_outs_15(scheduleDispatch_io_outs_15),
    .io_outs_14(scheduleDispatch_io_outs_14),
    .io_outs_13(scheduleDispatch_io_outs_13),
    .io_outs_12(scheduleDispatch_io_outs_12),
    .io_outs_11(scheduleDispatch_io_outs_11),
    .io_outs_10(scheduleDispatch_io_outs_10),
    .io_outs_9(scheduleDispatch_io_outs_9),
    .io_outs_8(scheduleDispatch_io_outs_8),
    .io_outs_7(scheduleDispatch_io_outs_7),
    .io_outs_6(scheduleDispatch_io_outs_6),
    .io_outs_5(scheduleDispatch_io_outs_5),
    .io_outs_4(scheduleDispatch_io_outs_4),
    .io_outs_3(scheduleDispatch_io_outs_3),
    .io_outs_2(scheduleDispatch_io_outs_2),
    .io_outs_1(scheduleDispatch_io_outs_1),
    .io_outs_0(scheduleDispatch_io_outs_0)
  );
  Alu Alu ( // @[TopModule.scala 124:54]
    .clock(Alu_clock),
    .reset(Alu_reset),
    .io_en(Alu_io_en),
    .io_skewing(Alu_io_skewing),
    .io_configuration(Alu_io_configuration),
    .io_inputs_1(Alu_io_inputs_1),
    .io_inputs_0(Alu_io_inputs_0),
    .io_outs_0(Alu_io_outs_0)
  );
  Alu Alu_1 ( // @[TopModule.scala 124:54]
    .clock(Alu_1_clock),
    .reset(Alu_1_reset),
    .io_en(Alu_1_io_en),
    .io_skewing(Alu_1_io_skewing),
    .io_configuration(Alu_1_io_configuration),
    .io_inputs_1(Alu_1_io_inputs_1),
    .io_inputs_0(Alu_1_io_inputs_0),
    .io_outs_0(Alu_1_io_outs_0)
  );
  Alu Alu_2 ( // @[TopModule.scala 124:54]
    .clock(Alu_2_clock),
    .reset(Alu_2_reset),
    .io_en(Alu_2_io_en),
    .io_skewing(Alu_2_io_skewing),
    .io_configuration(Alu_2_io_configuration),
    .io_inputs_1(Alu_2_io_inputs_1),
    .io_inputs_0(Alu_2_io_inputs_0),
    .io_outs_0(Alu_2_io_outs_0)
  );
  Alu Alu_3 ( // @[TopModule.scala 124:54]
    .clock(Alu_3_clock),
    .reset(Alu_3_reset),
    .io_en(Alu_3_io_en),
    .io_skewing(Alu_3_io_skewing),
    .io_configuration(Alu_3_io_configuration),
    .io_inputs_1(Alu_3_io_inputs_1),
    .io_inputs_0(Alu_3_io_inputs_0),
    .io_outs_0(Alu_3_io_outs_0)
  );
  Alu Alu_4 ( // @[TopModule.scala 124:54]
    .clock(Alu_4_clock),
    .reset(Alu_4_reset),
    .io_en(Alu_4_io_en),
    .io_skewing(Alu_4_io_skewing),
    .io_configuration(Alu_4_io_configuration),
    .io_inputs_1(Alu_4_io_inputs_1),
    .io_inputs_0(Alu_4_io_inputs_0),
    .io_outs_0(Alu_4_io_outs_0)
  );
  Alu Alu_5 ( // @[TopModule.scala 124:54]
    .clock(Alu_5_clock),
    .reset(Alu_5_reset),
    .io_en(Alu_5_io_en),
    .io_skewing(Alu_5_io_skewing),
    .io_configuration(Alu_5_io_configuration),
    .io_inputs_1(Alu_5_io_inputs_1),
    .io_inputs_0(Alu_5_io_inputs_0),
    .io_outs_0(Alu_5_io_outs_0)
  );
  Alu Alu_6 ( // @[TopModule.scala 124:54]
    .clock(Alu_6_clock),
    .reset(Alu_6_reset),
    .io_en(Alu_6_io_en),
    .io_skewing(Alu_6_io_skewing),
    .io_configuration(Alu_6_io_configuration),
    .io_inputs_1(Alu_6_io_inputs_1),
    .io_inputs_0(Alu_6_io_inputs_0),
    .io_outs_0(Alu_6_io_outs_0)
  );
  Alu Alu_7 ( // @[TopModule.scala 124:54]
    .clock(Alu_7_clock),
    .reset(Alu_7_reset),
    .io_en(Alu_7_io_en),
    .io_skewing(Alu_7_io_skewing),
    .io_configuration(Alu_7_io_configuration),
    .io_inputs_1(Alu_7_io_inputs_1),
    .io_inputs_0(Alu_7_io_inputs_0),
    .io_outs_0(Alu_7_io_outs_0)
  );
  Alu Alu_8 ( // @[TopModule.scala 124:54]
    .clock(Alu_8_clock),
    .reset(Alu_8_reset),
    .io_en(Alu_8_io_en),
    .io_skewing(Alu_8_io_skewing),
    .io_configuration(Alu_8_io_configuration),
    .io_inputs_1(Alu_8_io_inputs_1),
    .io_inputs_0(Alu_8_io_inputs_0),
    .io_outs_0(Alu_8_io_outs_0)
  );
  Alu Alu_9 ( // @[TopModule.scala 124:54]
    .clock(Alu_9_clock),
    .reset(Alu_9_reset),
    .io_en(Alu_9_io_en),
    .io_skewing(Alu_9_io_skewing),
    .io_configuration(Alu_9_io_configuration),
    .io_inputs_1(Alu_9_io_inputs_1),
    .io_inputs_0(Alu_9_io_inputs_0),
    .io_outs_0(Alu_9_io_outs_0)
  );
  Alu Alu_10 ( // @[TopModule.scala 124:54]
    .clock(Alu_10_clock),
    .reset(Alu_10_reset),
    .io_en(Alu_10_io_en),
    .io_skewing(Alu_10_io_skewing),
    .io_configuration(Alu_10_io_configuration),
    .io_inputs_1(Alu_10_io_inputs_1),
    .io_inputs_0(Alu_10_io_inputs_0),
    .io_outs_0(Alu_10_io_outs_0)
  );
  Alu Alu_11 ( // @[TopModule.scala 124:54]
    .clock(Alu_11_clock),
    .reset(Alu_11_reset),
    .io_en(Alu_11_io_en),
    .io_skewing(Alu_11_io_skewing),
    .io_configuration(Alu_11_io_configuration),
    .io_inputs_1(Alu_11_io_inputs_1),
    .io_inputs_0(Alu_11_io_inputs_0),
    .io_outs_0(Alu_11_io_outs_0)
  );
  Alu Alu_12 ( // @[TopModule.scala 124:54]
    .clock(Alu_12_clock),
    .reset(Alu_12_reset),
    .io_en(Alu_12_io_en),
    .io_skewing(Alu_12_io_skewing),
    .io_configuration(Alu_12_io_configuration),
    .io_inputs_1(Alu_12_io_inputs_1),
    .io_inputs_0(Alu_12_io_inputs_0),
    .io_outs_0(Alu_12_io_outs_0)
  );
  Alu Alu_13 ( // @[TopModule.scala 124:54]
    .clock(Alu_13_clock),
    .reset(Alu_13_reset),
    .io_en(Alu_13_io_en),
    .io_skewing(Alu_13_io_skewing),
    .io_configuration(Alu_13_io_configuration),
    .io_inputs_1(Alu_13_io_inputs_1),
    .io_inputs_0(Alu_13_io_inputs_0),
    .io_outs_0(Alu_13_io_outs_0)
  );
  Alu Alu_14 ( // @[TopModule.scala 124:54]
    .clock(Alu_14_clock),
    .reset(Alu_14_reset),
    .io_en(Alu_14_io_en),
    .io_skewing(Alu_14_io_skewing),
    .io_configuration(Alu_14_io_configuration),
    .io_inputs_1(Alu_14_io_inputs_1),
    .io_inputs_0(Alu_14_io_inputs_0),
    .io_outs_0(Alu_14_io_outs_0)
  );
  Alu Alu_15 ( // @[TopModule.scala 124:54]
    .clock(Alu_15_clock),
    .reset(Alu_15_reset),
    .io_en(Alu_15_io_en),
    .io_skewing(Alu_15_io_skewing),
    .io_configuration(Alu_15_io_configuration),
    .io_inputs_1(Alu_15_io_inputs_1),
    .io_inputs_0(Alu_15_io_inputs_0),
    .io_outs_0(Alu_15_io_outs_0)
  );
  MultiIIScheduleController MultiIIScheduleController ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_clock),
    .reset(MultiIIScheduleController_reset),
    .io_en(MultiIIScheduleController_io_en),
    .io_schedules_0(MultiIIScheduleController_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_io_schedules_3),
    .io_II(MultiIIScheduleController_io_II),
    .io_valid(MultiIIScheduleController_io_valid),
    .io_skewing(MultiIIScheduleController_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_1 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_1_clock),
    .reset(MultiIIScheduleController_1_reset),
    .io_en(MultiIIScheduleController_1_io_en),
    .io_schedules_0(MultiIIScheduleController_1_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_1_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_1_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_1_io_schedules_3),
    .io_II(MultiIIScheduleController_1_io_II),
    .io_valid(MultiIIScheduleController_1_io_valid),
    .io_skewing(MultiIIScheduleController_1_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_2 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_2_clock),
    .reset(MultiIIScheduleController_2_reset),
    .io_en(MultiIIScheduleController_2_io_en),
    .io_schedules_0(MultiIIScheduleController_2_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_2_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_2_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_2_io_schedules_3),
    .io_II(MultiIIScheduleController_2_io_II),
    .io_valid(MultiIIScheduleController_2_io_valid),
    .io_skewing(MultiIIScheduleController_2_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_3 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_3_clock),
    .reset(MultiIIScheduleController_3_reset),
    .io_en(MultiIIScheduleController_3_io_en),
    .io_schedules_0(MultiIIScheduleController_3_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_3_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_3_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_3_io_schedules_3),
    .io_II(MultiIIScheduleController_3_io_II),
    .io_valid(MultiIIScheduleController_3_io_valid),
    .io_skewing(MultiIIScheduleController_3_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_4 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_4_clock),
    .reset(MultiIIScheduleController_4_reset),
    .io_en(MultiIIScheduleController_4_io_en),
    .io_schedules_0(MultiIIScheduleController_4_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_4_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_4_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_4_io_schedules_3),
    .io_II(MultiIIScheduleController_4_io_II),
    .io_valid(MultiIIScheduleController_4_io_valid),
    .io_skewing(MultiIIScheduleController_4_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_5 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_5_clock),
    .reset(MultiIIScheduleController_5_reset),
    .io_en(MultiIIScheduleController_5_io_en),
    .io_schedules_0(MultiIIScheduleController_5_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_5_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_5_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_5_io_schedules_3),
    .io_II(MultiIIScheduleController_5_io_II),
    .io_valid(MultiIIScheduleController_5_io_valid),
    .io_skewing(MultiIIScheduleController_5_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_6 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_6_clock),
    .reset(MultiIIScheduleController_6_reset),
    .io_en(MultiIIScheduleController_6_io_en),
    .io_schedules_0(MultiIIScheduleController_6_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_6_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_6_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_6_io_schedules_3),
    .io_II(MultiIIScheduleController_6_io_II),
    .io_valid(MultiIIScheduleController_6_io_valid),
    .io_skewing(MultiIIScheduleController_6_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_7 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_7_clock),
    .reset(MultiIIScheduleController_7_reset),
    .io_en(MultiIIScheduleController_7_io_en),
    .io_schedules_0(MultiIIScheduleController_7_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_7_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_7_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_7_io_schedules_3),
    .io_II(MultiIIScheduleController_7_io_II),
    .io_valid(MultiIIScheduleController_7_io_valid),
    .io_skewing(MultiIIScheduleController_7_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_8 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_8_clock),
    .reset(MultiIIScheduleController_8_reset),
    .io_en(MultiIIScheduleController_8_io_en),
    .io_schedules_0(MultiIIScheduleController_8_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_8_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_8_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_8_io_schedules_3),
    .io_II(MultiIIScheduleController_8_io_II),
    .io_valid(MultiIIScheduleController_8_io_valid),
    .io_skewing(MultiIIScheduleController_8_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_9 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_9_clock),
    .reset(MultiIIScheduleController_9_reset),
    .io_en(MultiIIScheduleController_9_io_en),
    .io_schedules_0(MultiIIScheduleController_9_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_9_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_9_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_9_io_schedules_3),
    .io_II(MultiIIScheduleController_9_io_II),
    .io_valid(MultiIIScheduleController_9_io_valid),
    .io_skewing(MultiIIScheduleController_9_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_10 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_10_clock),
    .reset(MultiIIScheduleController_10_reset),
    .io_en(MultiIIScheduleController_10_io_en),
    .io_schedules_0(MultiIIScheduleController_10_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_10_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_10_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_10_io_schedules_3),
    .io_II(MultiIIScheduleController_10_io_II),
    .io_valid(MultiIIScheduleController_10_io_valid),
    .io_skewing(MultiIIScheduleController_10_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_11 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_11_clock),
    .reset(MultiIIScheduleController_11_reset),
    .io_en(MultiIIScheduleController_11_io_en),
    .io_schedules_0(MultiIIScheduleController_11_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_11_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_11_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_11_io_schedules_3),
    .io_II(MultiIIScheduleController_11_io_II),
    .io_valid(MultiIIScheduleController_11_io_valid),
    .io_skewing(MultiIIScheduleController_11_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_12 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_12_clock),
    .reset(MultiIIScheduleController_12_reset),
    .io_en(MultiIIScheduleController_12_io_en),
    .io_schedules_0(MultiIIScheduleController_12_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_12_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_12_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_12_io_schedules_3),
    .io_II(MultiIIScheduleController_12_io_II),
    .io_valid(MultiIIScheduleController_12_io_valid),
    .io_skewing(MultiIIScheduleController_12_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_13 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_13_clock),
    .reset(MultiIIScheduleController_13_reset),
    .io_en(MultiIIScheduleController_13_io_en),
    .io_schedules_0(MultiIIScheduleController_13_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_13_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_13_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_13_io_schedules_3),
    .io_II(MultiIIScheduleController_13_io_II),
    .io_valid(MultiIIScheduleController_13_io_valid),
    .io_skewing(MultiIIScheduleController_13_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_14 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_14_clock),
    .reset(MultiIIScheduleController_14_reset),
    .io_en(MultiIIScheduleController_14_io_en),
    .io_schedules_0(MultiIIScheduleController_14_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_14_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_14_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_14_io_schedules_3),
    .io_II(MultiIIScheduleController_14_io_II),
    .io_valid(MultiIIScheduleController_14_io_valid),
    .io_skewing(MultiIIScheduleController_14_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_15 ( // @[TopModule.scala 126:72]
    .clock(MultiIIScheduleController_15_clock),
    .reset(MultiIIScheduleController_15_reset),
    .io_en(MultiIIScheduleController_15_io_en),
    .io_schedules_0(MultiIIScheduleController_15_io_schedules_0),
    .io_schedules_1(MultiIIScheduleController_15_io_schedules_1),
    .io_schedules_2(MultiIIScheduleController_15_io_schedules_2),
    .io_schedules_3(MultiIIScheduleController_15_io_schedules_3),
    .io_II(MultiIIScheduleController_15_io_II),
    .io_valid(MultiIIScheduleController_15_io_valid),
    .io_skewing(MultiIIScheduleController_15_io_skewing)
  );
  RegisterFile RegisterFile ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_clock),
    .reset(RegisterFile_reset),
    .io_configuration(RegisterFile_io_configuration),
    .io_inputs_0(RegisterFile_io_inputs_0),
    .io_outs_1(RegisterFile_io_outs_1),
    .io_outs_0(RegisterFile_io_outs_0)
  );
  RegisterFile RegisterFile_1 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_1_clock),
    .reset(RegisterFile_1_reset),
    .io_configuration(RegisterFile_1_io_configuration),
    .io_inputs_0(RegisterFile_1_io_inputs_0),
    .io_outs_1(RegisterFile_1_io_outs_1),
    .io_outs_0(RegisterFile_1_io_outs_0)
  );
  RegisterFile RegisterFile_2 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_2_clock),
    .reset(RegisterFile_2_reset),
    .io_configuration(RegisterFile_2_io_configuration),
    .io_inputs_0(RegisterFile_2_io_inputs_0),
    .io_outs_1(RegisterFile_2_io_outs_1),
    .io_outs_0(RegisterFile_2_io_outs_0)
  );
  RegisterFile RegisterFile_3 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_3_clock),
    .reset(RegisterFile_3_reset),
    .io_configuration(RegisterFile_3_io_configuration),
    .io_inputs_0(RegisterFile_3_io_inputs_0),
    .io_outs_1(RegisterFile_3_io_outs_1),
    .io_outs_0(RegisterFile_3_io_outs_0)
  );
  RegisterFile RegisterFile_4 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_4_clock),
    .reset(RegisterFile_4_reset),
    .io_configuration(RegisterFile_4_io_configuration),
    .io_inputs_0(RegisterFile_4_io_inputs_0),
    .io_outs_1(RegisterFile_4_io_outs_1),
    .io_outs_0(RegisterFile_4_io_outs_0)
  );
  RegisterFile RegisterFile_5 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_5_clock),
    .reset(RegisterFile_5_reset),
    .io_configuration(RegisterFile_5_io_configuration),
    .io_inputs_0(RegisterFile_5_io_inputs_0),
    .io_outs_1(RegisterFile_5_io_outs_1),
    .io_outs_0(RegisterFile_5_io_outs_0)
  );
  RegisterFile RegisterFile_6 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_6_clock),
    .reset(RegisterFile_6_reset),
    .io_configuration(RegisterFile_6_io_configuration),
    .io_inputs_0(RegisterFile_6_io_inputs_0),
    .io_outs_1(RegisterFile_6_io_outs_1),
    .io_outs_0(RegisterFile_6_io_outs_0)
  );
  RegisterFile RegisterFile_7 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_7_clock),
    .reset(RegisterFile_7_reset),
    .io_configuration(RegisterFile_7_io_configuration),
    .io_inputs_0(RegisterFile_7_io_inputs_0),
    .io_outs_1(RegisterFile_7_io_outs_1),
    .io_outs_0(RegisterFile_7_io_outs_0)
  );
  RegisterFile RegisterFile_8 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_8_clock),
    .reset(RegisterFile_8_reset),
    .io_configuration(RegisterFile_8_io_configuration),
    .io_inputs_0(RegisterFile_8_io_inputs_0),
    .io_outs_1(RegisterFile_8_io_outs_1),
    .io_outs_0(RegisterFile_8_io_outs_0)
  );
  RegisterFile RegisterFile_9 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_9_clock),
    .reset(RegisterFile_9_reset),
    .io_configuration(RegisterFile_9_io_configuration),
    .io_inputs_0(RegisterFile_9_io_inputs_0),
    .io_outs_1(RegisterFile_9_io_outs_1),
    .io_outs_0(RegisterFile_9_io_outs_0)
  );
  RegisterFile RegisterFile_10 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_10_clock),
    .reset(RegisterFile_10_reset),
    .io_configuration(RegisterFile_10_io_configuration),
    .io_inputs_0(RegisterFile_10_io_inputs_0),
    .io_outs_1(RegisterFile_10_io_outs_1),
    .io_outs_0(RegisterFile_10_io_outs_0)
  );
  RegisterFile RegisterFile_11 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_11_clock),
    .reset(RegisterFile_11_reset),
    .io_configuration(RegisterFile_11_io_configuration),
    .io_inputs_0(RegisterFile_11_io_inputs_0),
    .io_outs_1(RegisterFile_11_io_outs_1),
    .io_outs_0(RegisterFile_11_io_outs_0)
  );
  RegisterFile RegisterFile_12 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_12_clock),
    .reset(RegisterFile_12_reset),
    .io_configuration(RegisterFile_12_io_configuration),
    .io_inputs_0(RegisterFile_12_io_inputs_0),
    .io_outs_1(RegisterFile_12_io_outs_1),
    .io_outs_0(RegisterFile_12_io_outs_0)
  );
  RegisterFile RegisterFile_13 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_13_clock),
    .reset(RegisterFile_13_reset),
    .io_configuration(RegisterFile_13_io_configuration),
    .io_inputs_0(RegisterFile_13_io_inputs_0),
    .io_outs_1(RegisterFile_13_io_outs_1),
    .io_outs_0(RegisterFile_13_io_outs_0)
  );
  RegisterFile RegisterFile_14 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_14_clock),
    .reset(RegisterFile_14_reset),
    .io_configuration(RegisterFile_14_io_configuration),
    .io_inputs_0(RegisterFile_14_io_inputs_0),
    .io_outs_1(RegisterFile_14_io_outs_1),
    .io_outs_0(RegisterFile_14_io_outs_0)
  );
  RegisterFile RegisterFile_15 ( // @[TopModule.scala 142:21]
    .clock(RegisterFile_15_clock),
    .reset(RegisterFile_15_reset),
    .io_configuration(RegisterFile_15_io_configuration),
    .io_inputs_0(RegisterFile_15_io_inputs_0),
    .io_outs_1(RegisterFile_15_io_outs_1),
    .io_outs_0(RegisterFile_15_io_outs_0)
  );
  Multiplexer Multiplexer ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_io_configuration),
    .io_inputs_3(Multiplexer_io_inputs_3),
    .io_inputs_2(Multiplexer_io_inputs_2),
    .io_inputs_1(Multiplexer_io_inputs_1),
    .io_inputs_0(Multiplexer_io_inputs_0),
    .io_outs_0(Multiplexer_io_outs_0)
  );
  Multiplexer_1 Multiplexer_1 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_1_io_configuration),
    .io_inputs_1(Multiplexer_1_io_inputs_1),
    .io_inputs_0(Multiplexer_1_io_inputs_0),
    .io_outs_0(Multiplexer_1_io_outs_0)
  );
  Multiplexer_1 Multiplexer_2 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_2_io_configuration),
    .io_inputs_1(Multiplexer_2_io_inputs_1),
    .io_inputs_0(Multiplexer_2_io_inputs_0),
    .io_outs_0(Multiplexer_2_io_outs_0)
  );
  Multiplexer_1 Multiplexer_3 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_3_io_configuration),
    .io_inputs_1(Multiplexer_3_io_inputs_1),
    .io_inputs_0(Multiplexer_3_io_inputs_0),
    .io_outs_0(Multiplexer_3_io_outs_0)
  );
  Multiplexer_1 Multiplexer_4 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_4_io_configuration),
    .io_inputs_1(Multiplexer_4_io_inputs_1),
    .io_inputs_0(Multiplexer_4_io_inputs_0),
    .io_outs_0(Multiplexer_4_io_outs_0)
  );
  Multiplexer_5 Multiplexer_5 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_5_io_configuration),
    .io_inputs_5(Multiplexer_5_io_inputs_5),
    .io_inputs_4(Multiplexer_5_io_inputs_4),
    .io_inputs_3(Multiplexer_5_io_inputs_3),
    .io_inputs_2(Multiplexer_5_io_inputs_2),
    .io_inputs_1(Multiplexer_5_io_inputs_1),
    .io_inputs_0(Multiplexer_5_io_inputs_0),
    .io_outs_0(Multiplexer_5_io_outs_0)
  );
  Multiplexer_6 Multiplexer_6 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_6_io_configuration),
    .io_inputs_4(Multiplexer_6_io_inputs_4),
    .io_inputs_3(Multiplexer_6_io_inputs_3),
    .io_inputs_2(Multiplexer_6_io_inputs_2),
    .io_inputs_1(Multiplexer_6_io_inputs_1),
    .io_inputs_0(Multiplexer_6_io_inputs_0),
    .io_outs_0(Multiplexer_6_io_outs_0)
  );
  Multiplexer Multiplexer_7 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_7_io_configuration),
    .io_inputs_3(Multiplexer_7_io_inputs_3),
    .io_inputs_2(Multiplexer_7_io_inputs_2),
    .io_inputs_1(Multiplexer_7_io_inputs_1),
    .io_inputs_0(Multiplexer_7_io_inputs_0),
    .io_outs_0(Multiplexer_7_io_outs_0)
  );
  Multiplexer_1 Multiplexer_8 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_8_io_configuration),
    .io_inputs_1(Multiplexer_8_io_inputs_1),
    .io_inputs_0(Multiplexer_8_io_inputs_0),
    .io_outs_0(Multiplexer_8_io_outs_0)
  );
  Multiplexer_5 Multiplexer_9 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_9_io_configuration),
    .io_inputs_5(Multiplexer_9_io_inputs_5),
    .io_inputs_4(Multiplexer_9_io_inputs_4),
    .io_inputs_3(Multiplexer_9_io_inputs_3),
    .io_inputs_2(Multiplexer_9_io_inputs_2),
    .io_inputs_1(Multiplexer_9_io_inputs_1),
    .io_inputs_0(Multiplexer_9_io_inputs_0),
    .io_outs_0(Multiplexer_9_io_outs_0)
  );
  Multiplexer_6 Multiplexer_10 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_10_io_configuration),
    .io_inputs_4(Multiplexer_10_io_inputs_4),
    .io_inputs_3(Multiplexer_10_io_inputs_3),
    .io_inputs_2(Multiplexer_10_io_inputs_2),
    .io_inputs_1(Multiplexer_10_io_inputs_1),
    .io_inputs_0(Multiplexer_10_io_inputs_0),
    .io_outs_0(Multiplexer_10_io_outs_0)
  );
  Multiplexer Multiplexer_11 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_11_io_configuration),
    .io_inputs_3(Multiplexer_11_io_inputs_3),
    .io_inputs_2(Multiplexer_11_io_inputs_2),
    .io_inputs_1(Multiplexer_11_io_inputs_1),
    .io_inputs_0(Multiplexer_11_io_inputs_0),
    .io_outs_0(Multiplexer_11_io_outs_0)
  );
  Multiplexer_1 Multiplexer_12 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_12_io_configuration),
    .io_inputs_1(Multiplexer_12_io_inputs_1),
    .io_inputs_0(Multiplexer_12_io_inputs_0),
    .io_outs_0(Multiplexer_12_io_outs_0)
  );
  Multiplexer_5 Multiplexer_13 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_13_io_configuration),
    .io_inputs_5(Multiplexer_13_io_inputs_5),
    .io_inputs_4(Multiplexer_13_io_inputs_4),
    .io_inputs_3(Multiplexer_13_io_inputs_3),
    .io_inputs_2(Multiplexer_13_io_inputs_2),
    .io_inputs_1(Multiplexer_13_io_inputs_1),
    .io_inputs_0(Multiplexer_13_io_inputs_0),
    .io_outs_0(Multiplexer_13_io_outs_0)
  );
  Multiplexer_6 Multiplexer_14 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_14_io_configuration),
    .io_inputs_4(Multiplexer_14_io_inputs_4),
    .io_inputs_3(Multiplexer_14_io_inputs_3),
    .io_inputs_2(Multiplexer_14_io_inputs_2),
    .io_inputs_1(Multiplexer_14_io_inputs_1),
    .io_inputs_0(Multiplexer_14_io_inputs_0),
    .io_outs_0(Multiplexer_14_io_outs_0)
  );
  Multiplexer Multiplexer_15 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_15_io_configuration),
    .io_inputs_3(Multiplexer_15_io_inputs_3),
    .io_inputs_2(Multiplexer_15_io_inputs_2),
    .io_inputs_1(Multiplexer_15_io_inputs_1),
    .io_inputs_0(Multiplexer_15_io_inputs_0),
    .io_outs_0(Multiplexer_15_io_outs_0)
  );
  Multiplexer_1 Multiplexer_16 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_16_io_configuration),
    .io_inputs_1(Multiplexer_16_io_inputs_1),
    .io_inputs_0(Multiplexer_16_io_inputs_0),
    .io_outs_0(Multiplexer_16_io_outs_0)
  );
  Multiplexer_5 Multiplexer_17 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_17_io_configuration),
    .io_inputs_5(Multiplexer_17_io_inputs_5),
    .io_inputs_4(Multiplexer_17_io_inputs_4),
    .io_inputs_3(Multiplexer_17_io_inputs_3),
    .io_inputs_2(Multiplexer_17_io_inputs_2),
    .io_inputs_1(Multiplexer_17_io_inputs_1),
    .io_inputs_0(Multiplexer_17_io_inputs_0),
    .io_outs_0(Multiplexer_17_io_outs_0)
  );
  Multiplexer_6 Multiplexer_18 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_18_io_configuration),
    .io_inputs_4(Multiplexer_18_io_inputs_4),
    .io_inputs_3(Multiplexer_18_io_inputs_3),
    .io_inputs_2(Multiplexer_18_io_inputs_2),
    .io_inputs_1(Multiplexer_18_io_inputs_1),
    .io_inputs_0(Multiplexer_18_io_inputs_0),
    .io_outs_0(Multiplexer_18_io_outs_0)
  );
  Multiplexer Multiplexer_19 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_19_io_configuration),
    .io_inputs_3(Multiplexer_19_io_inputs_3),
    .io_inputs_2(Multiplexer_19_io_inputs_2),
    .io_inputs_1(Multiplexer_19_io_inputs_1),
    .io_inputs_0(Multiplexer_19_io_inputs_0),
    .io_outs_0(Multiplexer_19_io_outs_0)
  );
  Multiplexer_1 Multiplexer_20 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_20_io_configuration),
    .io_inputs_1(Multiplexer_20_io_inputs_1),
    .io_inputs_0(Multiplexer_20_io_inputs_0),
    .io_outs_0(Multiplexer_20_io_outs_0)
  );
  Multiplexer_5 Multiplexer_21 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_21_io_configuration),
    .io_inputs_5(Multiplexer_21_io_inputs_5),
    .io_inputs_4(Multiplexer_21_io_inputs_4),
    .io_inputs_3(Multiplexer_21_io_inputs_3),
    .io_inputs_2(Multiplexer_21_io_inputs_2),
    .io_inputs_1(Multiplexer_21_io_inputs_1),
    .io_inputs_0(Multiplexer_21_io_inputs_0),
    .io_outs_0(Multiplexer_21_io_outs_0)
  );
  Multiplexer_6 Multiplexer_22 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_22_io_configuration),
    .io_inputs_4(Multiplexer_22_io_inputs_4),
    .io_inputs_3(Multiplexer_22_io_inputs_3),
    .io_inputs_2(Multiplexer_22_io_inputs_2),
    .io_inputs_1(Multiplexer_22_io_inputs_1),
    .io_inputs_0(Multiplexer_22_io_inputs_0),
    .io_outs_0(Multiplexer_22_io_outs_0)
  );
  Multiplexer Multiplexer_23 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_23_io_configuration),
    .io_inputs_3(Multiplexer_23_io_inputs_3),
    .io_inputs_2(Multiplexer_23_io_inputs_2),
    .io_inputs_1(Multiplexer_23_io_inputs_1),
    .io_inputs_0(Multiplexer_23_io_inputs_0),
    .io_outs_0(Multiplexer_23_io_outs_0)
  );
  Multiplexer_1 Multiplexer_24 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_24_io_configuration),
    .io_inputs_1(Multiplexer_24_io_inputs_1),
    .io_inputs_0(Multiplexer_24_io_inputs_0),
    .io_outs_0(Multiplexer_24_io_outs_0)
  );
  Multiplexer_5 Multiplexer_25 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_25_io_configuration),
    .io_inputs_5(Multiplexer_25_io_inputs_5),
    .io_inputs_4(Multiplexer_25_io_inputs_4),
    .io_inputs_3(Multiplexer_25_io_inputs_3),
    .io_inputs_2(Multiplexer_25_io_inputs_2),
    .io_inputs_1(Multiplexer_25_io_inputs_1),
    .io_inputs_0(Multiplexer_25_io_inputs_0),
    .io_outs_0(Multiplexer_25_io_outs_0)
  );
  Multiplexer_6 Multiplexer_26 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_26_io_configuration),
    .io_inputs_4(Multiplexer_26_io_inputs_4),
    .io_inputs_3(Multiplexer_26_io_inputs_3),
    .io_inputs_2(Multiplexer_26_io_inputs_2),
    .io_inputs_1(Multiplexer_26_io_inputs_1),
    .io_inputs_0(Multiplexer_26_io_inputs_0),
    .io_outs_0(Multiplexer_26_io_outs_0)
  );
  Multiplexer Multiplexer_27 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_27_io_configuration),
    .io_inputs_3(Multiplexer_27_io_inputs_3),
    .io_inputs_2(Multiplexer_27_io_inputs_2),
    .io_inputs_1(Multiplexer_27_io_inputs_1),
    .io_inputs_0(Multiplexer_27_io_inputs_0),
    .io_outs_0(Multiplexer_27_io_outs_0)
  );
  Multiplexer_1 Multiplexer_28 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_28_io_configuration),
    .io_inputs_1(Multiplexer_28_io_inputs_1),
    .io_inputs_0(Multiplexer_28_io_inputs_0),
    .io_outs_0(Multiplexer_28_io_outs_0)
  );
  Multiplexer_5 Multiplexer_29 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_29_io_configuration),
    .io_inputs_5(Multiplexer_29_io_inputs_5),
    .io_inputs_4(Multiplexer_29_io_inputs_4),
    .io_inputs_3(Multiplexer_29_io_inputs_3),
    .io_inputs_2(Multiplexer_29_io_inputs_2),
    .io_inputs_1(Multiplexer_29_io_inputs_1),
    .io_inputs_0(Multiplexer_29_io_inputs_0),
    .io_outs_0(Multiplexer_29_io_outs_0)
  );
  Multiplexer_6 Multiplexer_30 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_30_io_configuration),
    .io_inputs_4(Multiplexer_30_io_inputs_4),
    .io_inputs_3(Multiplexer_30_io_inputs_3),
    .io_inputs_2(Multiplexer_30_io_inputs_2),
    .io_inputs_1(Multiplexer_30_io_inputs_1),
    .io_inputs_0(Multiplexer_30_io_inputs_0),
    .io_outs_0(Multiplexer_30_io_outs_0)
  );
  Multiplexer Multiplexer_31 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_31_io_configuration),
    .io_inputs_3(Multiplexer_31_io_inputs_3),
    .io_inputs_2(Multiplexer_31_io_inputs_2),
    .io_inputs_1(Multiplexer_31_io_inputs_1),
    .io_inputs_0(Multiplexer_31_io_inputs_0),
    .io_outs_0(Multiplexer_31_io_outs_0)
  );
  Multiplexer_1 Multiplexer_32 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_32_io_configuration),
    .io_inputs_1(Multiplexer_32_io_inputs_1),
    .io_inputs_0(Multiplexer_32_io_inputs_0),
    .io_outs_0(Multiplexer_32_io_outs_0)
  );
  Multiplexer_5 Multiplexer_33 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_33_io_configuration),
    .io_inputs_5(Multiplexer_33_io_inputs_5),
    .io_inputs_4(Multiplexer_33_io_inputs_4),
    .io_inputs_3(Multiplexer_33_io_inputs_3),
    .io_inputs_2(Multiplexer_33_io_inputs_2),
    .io_inputs_1(Multiplexer_33_io_inputs_1),
    .io_inputs_0(Multiplexer_33_io_inputs_0),
    .io_outs_0(Multiplexer_33_io_outs_0)
  );
  Multiplexer_6 Multiplexer_34 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_34_io_configuration),
    .io_inputs_4(Multiplexer_34_io_inputs_4),
    .io_inputs_3(Multiplexer_34_io_inputs_3),
    .io_inputs_2(Multiplexer_34_io_inputs_2),
    .io_inputs_1(Multiplexer_34_io_inputs_1),
    .io_inputs_0(Multiplexer_34_io_inputs_0),
    .io_outs_0(Multiplexer_34_io_outs_0)
  );
  Multiplexer Multiplexer_35 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_35_io_configuration),
    .io_inputs_3(Multiplexer_35_io_inputs_3),
    .io_inputs_2(Multiplexer_35_io_inputs_2),
    .io_inputs_1(Multiplexer_35_io_inputs_1),
    .io_inputs_0(Multiplexer_35_io_inputs_0),
    .io_outs_0(Multiplexer_35_io_outs_0)
  );
  Multiplexer_1 Multiplexer_36 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_36_io_configuration),
    .io_inputs_1(Multiplexer_36_io_inputs_1),
    .io_inputs_0(Multiplexer_36_io_inputs_0),
    .io_outs_0(Multiplexer_36_io_outs_0)
  );
  Multiplexer_5 Multiplexer_37 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_37_io_configuration),
    .io_inputs_5(Multiplexer_37_io_inputs_5),
    .io_inputs_4(Multiplexer_37_io_inputs_4),
    .io_inputs_3(Multiplexer_37_io_inputs_3),
    .io_inputs_2(Multiplexer_37_io_inputs_2),
    .io_inputs_1(Multiplexer_37_io_inputs_1),
    .io_inputs_0(Multiplexer_37_io_inputs_0),
    .io_outs_0(Multiplexer_37_io_outs_0)
  );
  Multiplexer_6 Multiplexer_38 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_38_io_configuration),
    .io_inputs_4(Multiplexer_38_io_inputs_4),
    .io_inputs_3(Multiplexer_38_io_inputs_3),
    .io_inputs_2(Multiplexer_38_io_inputs_2),
    .io_inputs_1(Multiplexer_38_io_inputs_1),
    .io_inputs_0(Multiplexer_38_io_inputs_0),
    .io_outs_0(Multiplexer_38_io_outs_0)
  );
  Multiplexer Multiplexer_39 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_39_io_configuration),
    .io_inputs_3(Multiplexer_39_io_inputs_3),
    .io_inputs_2(Multiplexer_39_io_inputs_2),
    .io_inputs_1(Multiplexer_39_io_inputs_1),
    .io_inputs_0(Multiplexer_39_io_inputs_0),
    .io_outs_0(Multiplexer_39_io_outs_0)
  );
  Multiplexer_1 Multiplexer_40 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_40_io_configuration),
    .io_inputs_1(Multiplexer_40_io_inputs_1),
    .io_inputs_0(Multiplexer_40_io_inputs_0),
    .io_outs_0(Multiplexer_40_io_outs_0)
  );
  Multiplexer_5 Multiplexer_41 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_41_io_configuration),
    .io_inputs_5(Multiplexer_41_io_inputs_5),
    .io_inputs_4(Multiplexer_41_io_inputs_4),
    .io_inputs_3(Multiplexer_41_io_inputs_3),
    .io_inputs_2(Multiplexer_41_io_inputs_2),
    .io_inputs_1(Multiplexer_41_io_inputs_1),
    .io_inputs_0(Multiplexer_41_io_inputs_0),
    .io_outs_0(Multiplexer_41_io_outs_0)
  );
  Multiplexer_6 Multiplexer_42 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_42_io_configuration),
    .io_inputs_4(Multiplexer_42_io_inputs_4),
    .io_inputs_3(Multiplexer_42_io_inputs_3),
    .io_inputs_2(Multiplexer_42_io_inputs_2),
    .io_inputs_1(Multiplexer_42_io_inputs_1),
    .io_inputs_0(Multiplexer_42_io_inputs_0),
    .io_outs_0(Multiplexer_42_io_outs_0)
  );
  Multiplexer Multiplexer_43 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_43_io_configuration),
    .io_inputs_3(Multiplexer_43_io_inputs_3),
    .io_inputs_2(Multiplexer_43_io_inputs_2),
    .io_inputs_1(Multiplexer_43_io_inputs_1),
    .io_inputs_0(Multiplexer_43_io_inputs_0),
    .io_outs_0(Multiplexer_43_io_outs_0)
  );
  Multiplexer_1 Multiplexer_44 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_44_io_configuration),
    .io_inputs_1(Multiplexer_44_io_inputs_1),
    .io_inputs_0(Multiplexer_44_io_inputs_0),
    .io_outs_0(Multiplexer_44_io_outs_0)
  );
  Multiplexer_5 Multiplexer_45 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_45_io_configuration),
    .io_inputs_5(Multiplexer_45_io_inputs_5),
    .io_inputs_4(Multiplexer_45_io_inputs_4),
    .io_inputs_3(Multiplexer_45_io_inputs_3),
    .io_inputs_2(Multiplexer_45_io_inputs_2),
    .io_inputs_1(Multiplexer_45_io_inputs_1),
    .io_inputs_0(Multiplexer_45_io_inputs_0),
    .io_outs_0(Multiplexer_45_io_outs_0)
  );
  Multiplexer_6 Multiplexer_46 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_46_io_configuration),
    .io_inputs_4(Multiplexer_46_io_inputs_4),
    .io_inputs_3(Multiplexer_46_io_inputs_3),
    .io_inputs_2(Multiplexer_46_io_inputs_2),
    .io_inputs_1(Multiplexer_46_io_inputs_1),
    .io_inputs_0(Multiplexer_46_io_inputs_0),
    .io_outs_0(Multiplexer_46_io_outs_0)
  );
  Multiplexer Multiplexer_47 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_47_io_configuration),
    .io_inputs_3(Multiplexer_47_io_inputs_3),
    .io_inputs_2(Multiplexer_47_io_inputs_2),
    .io_inputs_1(Multiplexer_47_io_inputs_1),
    .io_inputs_0(Multiplexer_47_io_inputs_0),
    .io_outs_0(Multiplexer_47_io_outs_0)
  );
  Multiplexer_1 Multiplexer_48 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_48_io_configuration),
    .io_inputs_1(Multiplexer_48_io_inputs_1),
    .io_inputs_0(Multiplexer_48_io_inputs_0),
    .io_outs_0(Multiplexer_48_io_outs_0)
  );
  Multiplexer_5 Multiplexer_49 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_49_io_configuration),
    .io_inputs_5(Multiplexer_49_io_inputs_5),
    .io_inputs_4(Multiplexer_49_io_inputs_4),
    .io_inputs_3(Multiplexer_49_io_inputs_3),
    .io_inputs_2(Multiplexer_49_io_inputs_2),
    .io_inputs_1(Multiplexer_49_io_inputs_1),
    .io_inputs_0(Multiplexer_49_io_inputs_0),
    .io_outs_0(Multiplexer_49_io_outs_0)
  );
  Multiplexer_6 Multiplexer_50 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_50_io_configuration),
    .io_inputs_4(Multiplexer_50_io_inputs_4),
    .io_inputs_3(Multiplexer_50_io_inputs_3),
    .io_inputs_2(Multiplexer_50_io_inputs_2),
    .io_inputs_1(Multiplexer_50_io_inputs_1),
    .io_inputs_0(Multiplexer_50_io_inputs_0),
    .io_outs_0(Multiplexer_50_io_outs_0)
  );
  Multiplexer Multiplexer_51 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_51_io_configuration),
    .io_inputs_3(Multiplexer_51_io_inputs_3),
    .io_inputs_2(Multiplexer_51_io_inputs_2),
    .io_inputs_1(Multiplexer_51_io_inputs_1),
    .io_inputs_0(Multiplexer_51_io_inputs_0),
    .io_outs_0(Multiplexer_51_io_outs_0)
  );
  Multiplexer_1 Multiplexer_52 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_52_io_configuration),
    .io_inputs_1(Multiplexer_52_io_inputs_1),
    .io_inputs_0(Multiplexer_52_io_inputs_0),
    .io_outs_0(Multiplexer_52_io_outs_0)
  );
  Multiplexer_5 Multiplexer_53 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_53_io_configuration),
    .io_inputs_5(Multiplexer_53_io_inputs_5),
    .io_inputs_4(Multiplexer_53_io_inputs_4),
    .io_inputs_3(Multiplexer_53_io_inputs_3),
    .io_inputs_2(Multiplexer_53_io_inputs_2),
    .io_inputs_1(Multiplexer_53_io_inputs_1),
    .io_inputs_0(Multiplexer_53_io_inputs_0),
    .io_outs_0(Multiplexer_53_io_outs_0)
  );
  Multiplexer_6 Multiplexer_54 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_54_io_configuration),
    .io_inputs_4(Multiplexer_54_io_inputs_4),
    .io_inputs_3(Multiplexer_54_io_inputs_3),
    .io_inputs_2(Multiplexer_54_io_inputs_2),
    .io_inputs_1(Multiplexer_54_io_inputs_1),
    .io_inputs_0(Multiplexer_54_io_inputs_0),
    .io_outs_0(Multiplexer_54_io_outs_0)
  );
  Multiplexer Multiplexer_55 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_55_io_configuration),
    .io_inputs_3(Multiplexer_55_io_inputs_3),
    .io_inputs_2(Multiplexer_55_io_inputs_2),
    .io_inputs_1(Multiplexer_55_io_inputs_1),
    .io_inputs_0(Multiplexer_55_io_inputs_0),
    .io_outs_0(Multiplexer_55_io_outs_0)
  );
  Multiplexer_1 Multiplexer_56 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_56_io_configuration),
    .io_inputs_1(Multiplexer_56_io_inputs_1),
    .io_inputs_0(Multiplexer_56_io_inputs_0),
    .io_outs_0(Multiplexer_56_io_outs_0)
  );
  Multiplexer_5 Multiplexer_57 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_57_io_configuration),
    .io_inputs_5(Multiplexer_57_io_inputs_5),
    .io_inputs_4(Multiplexer_57_io_inputs_4),
    .io_inputs_3(Multiplexer_57_io_inputs_3),
    .io_inputs_2(Multiplexer_57_io_inputs_2),
    .io_inputs_1(Multiplexer_57_io_inputs_1),
    .io_inputs_0(Multiplexer_57_io_inputs_0),
    .io_outs_0(Multiplexer_57_io_outs_0)
  );
  Multiplexer_6 Multiplexer_58 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_58_io_configuration),
    .io_inputs_4(Multiplexer_58_io_inputs_4),
    .io_inputs_3(Multiplexer_58_io_inputs_3),
    .io_inputs_2(Multiplexer_58_io_inputs_2),
    .io_inputs_1(Multiplexer_58_io_inputs_1),
    .io_inputs_0(Multiplexer_58_io_inputs_0),
    .io_outs_0(Multiplexer_58_io_outs_0)
  );
  Multiplexer Multiplexer_59 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_59_io_configuration),
    .io_inputs_3(Multiplexer_59_io_inputs_3),
    .io_inputs_2(Multiplexer_59_io_inputs_2),
    .io_inputs_1(Multiplexer_59_io_inputs_1),
    .io_inputs_0(Multiplexer_59_io_inputs_0),
    .io_outs_0(Multiplexer_59_io_outs_0)
  );
  Multiplexer_1 Multiplexer_60 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_60_io_configuration),
    .io_inputs_1(Multiplexer_60_io_inputs_1),
    .io_inputs_0(Multiplexer_60_io_inputs_0),
    .io_outs_0(Multiplexer_60_io_outs_0)
  );
  Multiplexer_5 Multiplexer_61 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_61_io_configuration),
    .io_inputs_5(Multiplexer_61_io_inputs_5),
    .io_inputs_4(Multiplexer_61_io_inputs_4),
    .io_inputs_3(Multiplexer_61_io_inputs_3),
    .io_inputs_2(Multiplexer_61_io_inputs_2),
    .io_inputs_1(Multiplexer_61_io_inputs_1),
    .io_inputs_0(Multiplexer_61_io_inputs_0),
    .io_outs_0(Multiplexer_61_io_outs_0)
  );
  Multiplexer_6 Multiplexer_62 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_62_io_configuration),
    .io_inputs_4(Multiplexer_62_io_inputs_4),
    .io_inputs_3(Multiplexer_62_io_inputs_3),
    .io_inputs_2(Multiplexer_62_io_inputs_2),
    .io_inputs_1(Multiplexer_62_io_inputs_1),
    .io_inputs_0(Multiplexer_62_io_inputs_0),
    .io_outs_0(Multiplexer_62_io_outs_0)
  );
  Multiplexer Multiplexer_63 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_63_io_configuration),
    .io_inputs_3(Multiplexer_63_io_inputs_3),
    .io_inputs_2(Multiplexer_63_io_inputs_2),
    .io_inputs_1(Multiplexer_63_io_inputs_1),
    .io_inputs_0(Multiplexer_63_io_inputs_0),
    .io_outs_0(Multiplexer_63_io_outs_0)
  );
  Multiplexer_1 Multiplexer_64 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_64_io_configuration),
    .io_inputs_1(Multiplexer_64_io_inputs_1),
    .io_inputs_0(Multiplexer_64_io_inputs_0),
    .io_outs_0(Multiplexer_64_io_outs_0)
  );
  Multiplexer_5 Multiplexer_65 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_65_io_configuration),
    .io_inputs_5(Multiplexer_65_io_inputs_5),
    .io_inputs_4(Multiplexer_65_io_inputs_4),
    .io_inputs_3(Multiplexer_65_io_inputs_3),
    .io_inputs_2(Multiplexer_65_io_inputs_2),
    .io_inputs_1(Multiplexer_65_io_inputs_1),
    .io_inputs_0(Multiplexer_65_io_inputs_0),
    .io_outs_0(Multiplexer_65_io_outs_0)
  );
  Multiplexer_6 Multiplexer_66 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_66_io_configuration),
    .io_inputs_4(Multiplexer_66_io_inputs_4),
    .io_inputs_3(Multiplexer_66_io_inputs_3),
    .io_inputs_2(Multiplexer_66_io_inputs_2),
    .io_inputs_1(Multiplexer_66_io_inputs_1),
    .io_inputs_0(Multiplexer_66_io_inputs_0),
    .io_outs_0(Multiplexer_66_io_outs_0)
  );
  Multiplexer Multiplexer_67 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_67_io_configuration),
    .io_inputs_3(Multiplexer_67_io_inputs_3),
    .io_inputs_2(Multiplexer_67_io_inputs_2),
    .io_inputs_1(Multiplexer_67_io_inputs_1),
    .io_inputs_0(Multiplexer_67_io_inputs_0),
    .io_outs_0(Multiplexer_67_io_outs_0)
  );
  Multiplexer_1 Multiplexer_68 ( // @[TopModule.scala 153:11]
    .io_configuration(Multiplexer_68_io_configuration),
    .io_inputs_1(Multiplexer_68_io_inputs_1),
    .io_inputs_0(Multiplexer_68_io_inputs_0),
    .io_outs_0(Multiplexer_68_io_outs_0)
  );
  ConstUnit ConstUnit ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_io_configuration),
    .io_outs_0(ConstUnit_io_outs_0)
  );
  ConstUnit ConstUnit_1 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_1_io_configuration),
    .io_outs_0(ConstUnit_1_io_outs_0)
  );
  ConstUnit ConstUnit_2 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_2_io_configuration),
    .io_outs_0(ConstUnit_2_io_outs_0)
  );
  ConstUnit ConstUnit_3 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_3_io_configuration),
    .io_outs_0(ConstUnit_3_io_outs_0)
  );
  ConstUnit ConstUnit_4 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_4_io_configuration),
    .io_outs_0(ConstUnit_4_io_outs_0)
  );
  ConstUnit ConstUnit_5 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_5_io_configuration),
    .io_outs_0(ConstUnit_5_io_outs_0)
  );
  ConstUnit ConstUnit_6 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_6_io_configuration),
    .io_outs_0(ConstUnit_6_io_outs_0)
  );
  ConstUnit ConstUnit_7 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_7_io_configuration),
    .io_outs_0(ConstUnit_7_io_outs_0)
  );
  ConstUnit ConstUnit_8 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_8_io_configuration),
    .io_outs_0(ConstUnit_8_io_outs_0)
  );
  ConstUnit ConstUnit_9 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_9_io_configuration),
    .io_outs_0(ConstUnit_9_io_outs_0)
  );
  ConstUnit ConstUnit_10 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_10_io_configuration),
    .io_outs_0(ConstUnit_10_io_outs_0)
  );
  ConstUnit ConstUnit_11 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_11_io_configuration),
    .io_outs_0(ConstUnit_11_io_outs_0)
  );
  ConstUnit ConstUnit_12 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_12_io_configuration),
    .io_outs_0(ConstUnit_12_io_outs_0)
  );
  ConstUnit ConstUnit_13 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_13_io_configuration),
    .io_outs_0(ConstUnit_13_io_outs_0)
  );
  ConstUnit ConstUnit_14 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_14_io_configuration),
    .io_outs_0(ConstUnit_14_io_outs_0)
  );
  ConstUnit ConstUnit_15 ( // @[TopModule.scala 161:21]
    .io_configuration(ConstUnit_15_io_configuration),
    .io_outs_0(ConstUnit_15_io_outs_0)
  );
  ConfigController configControllers_0 ( // @[TopModule.scala 234:34]
    .clock(configControllers_0_clock),
    .reset(configControllers_0_reset),
    .io_en(configControllers_0_io_en),
    .io_II(configControllers_0_io_II),
    .io_inConfig(configControllers_0_io_inConfig),
    .io_outConfig(configControllers_0_io_outConfig)
  );
  Dispatch_17 Dispatch ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_io_configuration),
    .io_outs_4(Dispatch_io_outs_4),
    .io_outs_3(Dispatch_io_outs_3),
    .io_outs_2(Dispatch_io_outs_2),
    .io_outs_1(Dispatch_io_outs_1),
    .io_outs_0(Dispatch_io_outs_0)
  );
  ConfigController_1 configControllers_1 ( // @[TopModule.scala 234:34]
    .clock(configControllers_1_clock),
    .reset(configControllers_1_reset),
    .io_en(configControllers_1_io_en),
    .io_II(configControllers_1_io_II),
    .io_inConfig(configControllers_1_io_inConfig),
    .io_outConfig(configControllers_1_io_outConfig)
  );
  Dispatch_18 Dispatch_1 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_1_io_configuration),
    .io_outs_6(Dispatch_1_io_outs_6),
    .io_outs_5(Dispatch_1_io_outs_5),
    .io_outs_4(Dispatch_1_io_outs_4),
    .io_outs_3(Dispatch_1_io_outs_3),
    .io_outs_2(Dispatch_1_io_outs_2),
    .io_outs_1(Dispatch_1_io_outs_1),
    .io_outs_0(Dispatch_1_io_outs_0)
  );
  ConfigController_1 configControllers_2 ( // @[TopModule.scala 234:34]
    .clock(configControllers_2_clock),
    .reset(configControllers_2_reset),
    .io_en(configControllers_2_io_en),
    .io_II(configControllers_2_io_II),
    .io_inConfig(configControllers_2_io_inConfig),
    .io_outConfig(configControllers_2_io_outConfig)
  );
  Dispatch_18 Dispatch_2 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_2_io_configuration),
    .io_outs_6(Dispatch_2_io_outs_6),
    .io_outs_5(Dispatch_2_io_outs_5),
    .io_outs_4(Dispatch_2_io_outs_4),
    .io_outs_3(Dispatch_2_io_outs_3),
    .io_outs_2(Dispatch_2_io_outs_2),
    .io_outs_1(Dispatch_2_io_outs_1),
    .io_outs_0(Dispatch_2_io_outs_0)
  );
  ConfigController_1 configControllers_3 ( // @[TopModule.scala 234:34]
    .clock(configControllers_3_clock),
    .reset(configControllers_3_reset),
    .io_en(configControllers_3_io_en),
    .io_II(configControllers_3_io_II),
    .io_inConfig(configControllers_3_io_inConfig),
    .io_outConfig(configControllers_3_io_outConfig)
  );
  Dispatch_18 Dispatch_3 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_3_io_configuration),
    .io_outs_6(Dispatch_3_io_outs_6),
    .io_outs_5(Dispatch_3_io_outs_5),
    .io_outs_4(Dispatch_3_io_outs_4),
    .io_outs_3(Dispatch_3_io_outs_3),
    .io_outs_2(Dispatch_3_io_outs_2),
    .io_outs_1(Dispatch_3_io_outs_1),
    .io_outs_0(Dispatch_3_io_outs_0)
  );
  ConfigController_1 configControllers_4 ( // @[TopModule.scala 234:34]
    .clock(configControllers_4_clock),
    .reset(configControllers_4_reset),
    .io_en(configControllers_4_io_en),
    .io_II(configControllers_4_io_II),
    .io_inConfig(configControllers_4_io_inConfig),
    .io_outConfig(configControllers_4_io_outConfig)
  );
  Dispatch_18 Dispatch_4 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_4_io_configuration),
    .io_outs_6(Dispatch_4_io_outs_6),
    .io_outs_5(Dispatch_4_io_outs_5),
    .io_outs_4(Dispatch_4_io_outs_4),
    .io_outs_3(Dispatch_4_io_outs_3),
    .io_outs_2(Dispatch_4_io_outs_2),
    .io_outs_1(Dispatch_4_io_outs_1),
    .io_outs_0(Dispatch_4_io_outs_0)
  );
  ConfigController_1 configControllers_5 ( // @[TopModule.scala 234:34]
    .clock(configControllers_5_clock),
    .reset(configControllers_5_reset),
    .io_en(configControllers_5_io_en),
    .io_II(configControllers_5_io_II),
    .io_inConfig(configControllers_5_io_inConfig),
    .io_outConfig(configControllers_5_io_outConfig)
  );
  Dispatch_18 Dispatch_5 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_5_io_configuration),
    .io_outs_6(Dispatch_5_io_outs_6),
    .io_outs_5(Dispatch_5_io_outs_5),
    .io_outs_4(Dispatch_5_io_outs_4),
    .io_outs_3(Dispatch_5_io_outs_3),
    .io_outs_2(Dispatch_5_io_outs_2),
    .io_outs_1(Dispatch_5_io_outs_1),
    .io_outs_0(Dispatch_5_io_outs_0)
  );
  ConfigController_1 configControllers_6 ( // @[TopModule.scala 234:34]
    .clock(configControllers_6_clock),
    .reset(configControllers_6_reset),
    .io_en(configControllers_6_io_en),
    .io_II(configControllers_6_io_II),
    .io_inConfig(configControllers_6_io_inConfig),
    .io_outConfig(configControllers_6_io_outConfig)
  );
  Dispatch_18 Dispatch_6 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_6_io_configuration),
    .io_outs_6(Dispatch_6_io_outs_6),
    .io_outs_5(Dispatch_6_io_outs_5),
    .io_outs_4(Dispatch_6_io_outs_4),
    .io_outs_3(Dispatch_6_io_outs_3),
    .io_outs_2(Dispatch_6_io_outs_2),
    .io_outs_1(Dispatch_6_io_outs_1),
    .io_outs_0(Dispatch_6_io_outs_0)
  );
  ConfigController_1 configControllers_7 ( // @[TopModule.scala 234:34]
    .clock(configControllers_7_clock),
    .reset(configControllers_7_reset),
    .io_en(configControllers_7_io_en),
    .io_II(configControllers_7_io_II),
    .io_inConfig(configControllers_7_io_inConfig),
    .io_outConfig(configControllers_7_io_outConfig)
  );
  Dispatch_18 Dispatch_7 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_7_io_configuration),
    .io_outs_6(Dispatch_7_io_outs_6),
    .io_outs_5(Dispatch_7_io_outs_5),
    .io_outs_4(Dispatch_7_io_outs_4),
    .io_outs_3(Dispatch_7_io_outs_3),
    .io_outs_2(Dispatch_7_io_outs_2),
    .io_outs_1(Dispatch_7_io_outs_1),
    .io_outs_0(Dispatch_7_io_outs_0)
  );
  ConfigController_1 configControllers_8 ( // @[TopModule.scala 234:34]
    .clock(configControllers_8_clock),
    .reset(configControllers_8_reset),
    .io_en(configControllers_8_io_en),
    .io_II(configControllers_8_io_II),
    .io_inConfig(configControllers_8_io_inConfig),
    .io_outConfig(configControllers_8_io_outConfig)
  );
  Dispatch_18 Dispatch_8 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_8_io_configuration),
    .io_outs_6(Dispatch_8_io_outs_6),
    .io_outs_5(Dispatch_8_io_outs_5),
    .io_outs_4(Dispatch_8_io_outs_4),
    .io_outs_3(Dispatch_8_io_outs_3),
    .io_outs_2(Dispatch_8_io_outs_2),
    .io_outs_1(Dispatch_8_io_outs_1),
    .io_outs_0(Dispatch_8_io_outs_0)
  );
  ConfigController_1 configControllers_9 ( // @[TopModule.scala 234:34]
    .clock(configControllers_9_clock),
    .reset(configControllers_9_reset),
    .io_en(configControllers_9_io_en),
    .io_II(configControllers_9_io_II),
    .io_inConfig(configControllers_9_io_inConfig),
    .io_outConfig(configControllers_9_io_outConfig)
  );
  Dispatch_18 Dispatch_9 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_9_io_configuration),
    .io_outs_6(Dispatch_9_io_outs_6),
    .io_outs_5(Dispatch_9_io_outs_5),
    .io_outs_4(Dispatch_9_io_outs_4),
    .io_outs_3(Dispatch_9_io_outs_3),
    .io_outs_2(Dispatch_9_io_outs_2),
    .io_outs_1(Dispatch_9_io_outs_1),
    .io_outs_0(Dispatch_9_io_outs_0)
  );
  ConfigController_1 configControllers_10 ( // @[TopModule.scala 234:34]
    .clock(configControllers_10_clock),
    .reset(configControllers_10_reset),
    .io_en(configControllers_10_io_en),
    .io_II(configControllers_10_io_II),
    .io_inConfig(configControllers_10_io_inConfig),
    .io_outConfig(configControllers_10_io_outConfig)
  );
  Dispatch_18 Dispatch_10 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_10_io_configuration),
    .io_outs_6(Dispatch_10_io_outs_6),
    .io_outs_5(Dispatch_10_io_outs_5),
    .io_outs_4(Dispatch_10_io_outs_4),
    .io_outs_3(Dispatch_10_io_outs_3),
    .io_outs_2(Dispatch_10_io_outs_2),
    .io_outs_1(Dispatch_10_io_outs_1),
    .io_outs_0(Dispatch_10_io_outs_0)
  );
  ConfigController_1 configControllers_11 ( // @[TopModule.scala 234:34]
    .clock(configControllers_11_clock),
    .reset(configControllers_11_reset),
    .io_en(configControllers_11_io_en),
    .io_II(configControllers_11_io_II),
    .io_inConfig(configControllers_11_io_inConfig),
    .io_outConfig(configControllers_11_io_outConfig)
  );
  Dispatch_18 Dispatch_11 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_11_io_configuration),
    .io_outs_6(Dispatch_11_io_outs_6),
    .io_outs_5(Dispatch_11_io_outs_5),
    .io_outs_4(Dispatch_11_io_outs_4),
    .io_outs_3(Dispatch_11_io_outs_3),
    .io_outs_2(Dispatch_11_io_outs_2),
    .io_outs_1(Dispatch_11_io_outs_1),
    .io_outs_0(Dispatch_11_io_outs_0)
  );
  ConfigController_1 configControllers_12 ( // @[TopModule.scala 234:34]
    .clock(configControllers_12_clock),
    .reset(configControllers_12_reset),
    .io_en(configControllers_12_io_en),
    .io_II(configControllers_12_io_II),
    .io_inConfig(configControllers_12_io_inConfig),
    .io_outConfig(configControllers_12_io_outConfig)
  );
  Dispatch_18 Dispatch_12 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_12_io_configuration),
    .io_outs_6(Dispatch_12_io_outs_6),
    .io_outs_5(Dispatch_12_io_outs_5),
    .io_outs_4(Dispatch_12_io_outs_4),
    .io_outs_3(Dispatch_12_io_outs_3),
    .io_outs_2(Dispatch_12_io_outs_2),
    .io_outs_1(Dispatch_12_io_outs_1),
    .io_outs_0(Dispatch_12_io_outs_0)
  );
  ConfigController_1 configControllers_13 ( // @[TopModule.scala 234:34]
    .clock(configControllers_13_clock),
    .reset(configControllers_13_reset),
    .io_en(configControllers_13_io_en),
    .io_II(configControllers_13_io_II),
    .io_inConfig(configControllers_13_io_inConfig),
    .io_outConfig(configControllers_13_io_outConfig)
  );
  Dispatch_18 Dispatch_13 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_13_io_configuration),
    .io_outs_6(Dispatch_13_io_outs_6),
    .io_outs_5(Dispatch_13_io_outs_5),
    .io_outs_4(Dispatch_13_io_outs_4),
    .io_outs_3(Dispatch_13_io_outs_3),
    .io_outs_2(Dispatch_13_io_outs_2),
    .io_outs_1(Dispatch_13_io_outs_1),
    .io_outs_0(Dispatch_13_io_outs_0)
  );
  ConfigController_1 configControllers_14 ( // @[TopModule.scala 234:34]
    .clock(configControllers_14_clock),
    .reset(configControllers_14_reset),
    .io_en(configControllers_14_io_en),
    .io_II(configControllers_14_io_II),
    .io_inConfig(configControllers_14_io_inConfig),
    .io_outConfig(configControllers_14_io_outConfig)
  );
  Dispatch_18 Dispatch_14 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_14_io_configuration),
    .io_outs_6(Dispatch_14_io_outs_6),
    .io_outs_5(Dispatch_14_io_outs_5),
    .io_outs_4(Dispatch_14_io_outs_4),
    .io_outs_3(Dispatch_14_io_outs_3),
    .io_outs_2(Dispatch_14_io_outs_2),
    .io_outs_1(Dispatch_14_io_outs_1),
    .io_outs_0(Dispatch_14_io_outs_0)
  );
  ConfigController_1 configControllers_15 ( // @[TopModule.scala 234:34]
    .clock(configControllers_15_clock),
    .reset(configControllers_15_reset),
    .io_en(configControllers_15_io_en),
    .io_II(configControllers_15_io_II),
    .io_inConfig(configControllers_15_io_inConfig),
    .io_outConfig(configControllers_15_io_outConfig)
  );
  Dispatch_18 Dispatch_15 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_15_io_configuration),
    .io_outs_6(Dispatch_15_io_outs_6),
    .io_outs_5(Dispatch_15_io_outs_5),
    .io_outs_4(Dispatch_15_io_outs_4),
    .io_outs_3(Dispatch_15_io_outs_3),
    .io_outs_2(Dispatch_15_io_outs_2),
    .io_outs_1(Dispatch_15_io_outs_1),
    .io_outs_0(Dispatch_15_io_outs_0)
  );
  ConfigController_1 configControllers_16 ( // @[TopModule.scala 234:34]
    .clock(configControllers_16_clock),
    .reset(configControllers_16_reset),
    .io_en(configControllers_16_io_en),
    .io_II(configControllers_16_io_II),
    .io_inConfig(configControllers_16_io_inConfig),
    .io_outConfig(configControllers_16_io_outConfig)
  );
  Dispatch_18 Dispatch_16 ( // @[TopModule.scala 239:26]
    .io_configuration(Dispatch_16_io_configuration),
    .io_outs_6(Dispatch_16_io_outs_6),
    .io_outs_5(Dispatch_16_io_outs_5),
    .io_outs_4(Dispatch_16_io_outs_4),
    .io_outs_3(Dispatch_16_io_outs_3),
    .io_outs_2(Dispatch_16_io_outs_2),
    .io_outs_1(Dispatch_16_io_outs_1),
    .io_outs_0(Dispatch_16_io_outs_0)
  );
  Dispatch_34 topDispatch ( // @[TopModule.scala 248:27]
    .io_configuration(topDispatch_io_configuration),
    .io_outs_16(topDispatch_io_outs_16),
    .io_outs_15(topDispatch_io_outs_15),
    .io_outs_14(topDispatch_io_outs_14),
    .io_outs_13(topDispatch_io_outs_13),
    .io_outs_12(topDispatch_io_outs_12),
    .io_outs_11(topDispatch_io_outs_11),
    .io_outs_10(topDispatch_io_outs_10),
    .io_outs_9(topDispatch_io_outs_9),
    .io_outs_8(topDispatch_io_outs_8),
    .io_outs_7(topDispatch_io_outs_7),
    .io_outs_6(topDispatch_io_outs_6),
    .io_outs_5(topDispatch_io_outs_5),
    .io_outs_4(topDispatch_io_outs_4),
    .io_outs_3(topDispatch_io_outs_3),
    .io_outs_2(topDispatch_io_outs_2),
    .io_outs_1(topDispatch_io_outs_1),
    .io_outs_0(topDispatch_io_outs_0)
  );
  assign io_outs_0 = Multiplexer_io_outs_0; // @[TopModule.scala 263:25]
  assign scheduleDispatch_io_configuration = io_schedules; // @[TopModule.scala 120:37]
  assign Alu_clock = clock;
  assign Alu_reset = reset;
  assign Alu_io_en = MultiIIScheduleController_io_valid; // @[TopModule.scala 135:15]
  assign Alu_io_skewing = MultiIIScheduleController_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_io_configuration = Dispatch_1_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_io_inputs_1 = Multiplexer_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_io_inputs_0 = Multiplexer_5_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_1_clock = clock;
  assign Alu_1_reset = reset;
  assign Alu_1_io_en = MultiIIScheduleController_1_io_valid; // @[TopModule.scala 135:15]
  assign Alu_1_io_skewing = MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_1_io_configuration = Dispatch_2_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_1_io_inputs_1 = Multiplexer_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_1_io_inputs_0 = Multiplexer_9_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_2_clock = clock;
  assign Alu_2_reset = reset;
  assign Alu_2_io_en = MultiIIScheduleController_2_io_valid; // @[TopModule.scala 135:15]
  assign Alu_2_io_skewing = MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_2_io_configuration = Dispatch_3_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_2_io_inputs_1 = Multiplexer_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_2_io_inputs_0 = Multiplexer_13_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_3_clock = clock;
  assign Alu_3_reset = reset;
  assign Alu_3_io_en = MultiIIScheduleController_3_io_valid; // @[TopModule.scala 135:15]
  assign Alu_3_io_skewing = MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_3_io_configuration = Dispatch_4_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_3_io_inputs_1 = Multiplexer_18_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_3_io_inputs_0 = Multiplexer_17_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_4_clock = clock;
  assign Alu_4_reset = reset;
  assign Alu_4_io_en = MultiIIScheduleController_4_io_valid; // @[TopModule.scala 135:15]
  assign Alu_4_io_skewing = MultiIIScheduleController_4_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_4_io_configuration = Dispatch_5_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_4_io_inputs_1 = Multiplexer_22_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_4_io_inputs_0 = Multiplexer_21_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_5_clock = clock;
  assign Alu_5_reset = reset;
  assign Alu_5_io_en = MultiIIScheduleController_5_io_valid; // @[TopModule.scala 135:15]
  assign Alu_5_io_skewing = MultiIIScheduleController_5_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_5_io_configuration = Dispatch_6_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_5_io_inputs_1 = Multiplexer_26_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_5_io_inputs_0 = Multiplexer_25_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_6_clock = clock;
  assign Alu_6_reset = reset;
  assign Alu_6_io_en = MultiIIScheduleController_6_io_valid; // @[TopModule.scala 135:15]
  assign Alu_6_io_skewing = MultiIIScheduleController_6_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_6_io_configuration = Dispatch_7_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_6_io_inputs_1 = Multiplexer_30_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_6_io_inputs_0 = Multiplexer_29_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_7_clock = clock;
  assign Alu_7_reset = reset;
  assign Alu_7_io_en = MultiIIScheduleController_7_io_valid; // @[TopModule.scala 135:15]
  assign Alu_7_io_skewing = MultiIIScheduleController_7_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_7_io_configuration = Dispatch_8_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_7_io_inputs_1 = Multiplexer_34_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_7_io_inputs_0 = Multiplexer_33_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_8_clock = clock;
  assign Alu_8_reset = reset;
  assign Alu_8_io_en = MultiIIScheduleController_8_io_valid; // @[TopModule.scala 135:15]
  assign Alu_8_io_skewing = MultiIIScheduleController_8_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_8_io_configuration = Dispatch_9_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_8_io_inputs_1 = Multiplexer_38_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_8_io_inputs_0 = Multiplexer_37_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_9_clock = clock;
  assign Alu_9_reset = reset;
  assign Alu_9_io_en = MultiIIScheduleController_9_io_valid; // @[TopModule.scala 135:15]
  assign Alu_9_io_skewing = MultiIIScheduleController_9_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_9_io_configuration = Dispatch_10_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_9_io_inputs_1 = Multiplexer_42_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_9_io_inputs_0 = Multiplexer_41_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_10_clock = clock;
  assign Alu_10_reset = reset;
  assign Alu_10_io_en = MultiIIScheduleController_10_io_valid; // @[TopModule.scala 135:15]
  assign Alu_10_io_skewing = MultiIIScheduleController_10_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_10_io_configuration = Dispatch_11_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_10_io_inputs_1 = Multiplexer_46_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_10_io_inputs_0 = Multiplexer_45_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_11_clock = clock;
  assign Alu_11_reset = reset;
  assign Alu_11_io_en = MultiIIScheduleController_11_io_valid; // @[TopModule.scala 135:15]
  assign Alu_11_io_skewing = MultiIIScheduleController_11_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_11_io_configuration = Dispatch_12_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_11_io_inputs_1 = Multiplexer_50_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_11_io_inputs_0 = Multiplexer_49_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_12_clock = clock;
  assign Alu_12_reset = reset;
  assign Alu_12_io_en = MultiIIScheduleController_12_io_valid; // @[TopModule.scala 135:15]
  assign Alu_12_io_skewing = MultiIIScheduleController_12_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_12_io_configuration = Dispatch_13_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_12_io_inputs_1 = Multiplexer_54_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_12_io_inputs_0 = Multiplexer_53_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_13_clock = clock;
  assign Alu_13_reset = reset;
  assign Alu_13_io_en = MultiIIScheduleController_13_io_valid; // @[TopModule.scala 135:15]
  assign Alu_13_io_skewing = MultiIIScheduleController_13_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_13_io_configuration = Dispatch_14_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_13_io_inputs_1 = Multiplexer_58_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_13_io_inputs_0 = Multiplexer_57_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_14_clock = clock;
  assign Alu_14_reset = reset;
  assign Alu_14_io_en = MultiIIScheduleController_14_io_valid; // @[TopModule.scala 135:15]
  assign Alu_14_io_skewing = MultiIIScheduleController_14_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_14_io_configuration = Dispatch_15_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_14_io_inputs_1 = Multiplexer_62_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_14_io_inputs_0 = Multiplexer_61_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_15_clock = clock;
  assign Alu_15_reset = reset;
  assign Alu_15_io_en = MultiIIScheduleController_15_io_valid; // @[TopModule.scala 135:15]
  assign Alu_15_io_skewing = MultiIIScheduleController_15_io_skewing; // @[TopModule.scala 136:20]
  assign Alu_15_io_configuration = Dispatch_16_io_outs_0; // @[TopModule.scala 242:22]
  assign Alu_15_io_inputs_1 = Multiplexer_66_io_outs_0; // @[TopModule.scala 267:60]
  assign Alu_15_io_inputs_0 = Multiplexer_65_io_outs_0; // @[TopModule.scala 267:60]
  assign MultiIIScheduleController_clock = clock;
  assign MultiIIScheduleController_reset = reset;
  assign MultiIIScheduleController_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_io_schedules_0 = scheduleDispatch_io_outs_0; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_schedules_1 = scheduleDispatch_io_outs_1; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_schedules_2 = scheduleDispatch_io_outs_2; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_schedules_3 = scheduleDispatch_io_outs_3; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_1_clock = clock;
  assign MultiIIScheduleController_1_reset = reset;
  assign MultiIIScheduleController_1_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_1_io_schedules_0 = scheduleDispatch_io_outs_4; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_schedules_1 = scheduleDispatch_io_outs_5; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_schedules_2 = scheduleDispatch_io_outs_6; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_schedules_3 = scheduleDispatch_io_outs_7; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_1_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_2_clock = clock;
  assign MultiIIScheduleController_2_reset = reset;
  assign MultiIIScheduleController_2_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_2_io_schedules_0 = scheduleDispatch_io_outs_8; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_schedules_1 = scheduleDispatch_io_outs_9; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_schedules_2 = scheduleDispatch_io_outs_10; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_schedules_3 = scheduleDispatch_io_outs_11; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_2_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_3_clock = clock;
  assign MultiIIScheduleController_3_reset = reset;
  assign MultiIIScheduleController_3_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_3_io_schedules_0 = scheduleDispatch_io_outs_12; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_schedules_1 = scheduleDispatch_io_outs_13; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_schedules_2 = scheduleDispatch_io_outs_14; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_schedules_3 = scheduleDispatch_io_outs_15; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_3_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_4_clock = clock;
  assign MultiIIScheduleController_4_reset = reset;
  assign MultiIIScheduleController_4_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_4_io_schedules_0 = scheduleDispatch_io_outs_16; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_4_io_schedules_1 = scheduleDispatch_io_outs_17; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_4_io_schedules_2 = scheduleDispatch_io_outs_18; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_4_io_schedules_3 = scheduleDispatch_io_outs_19; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_4_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_5_clock = clock;
  assign MultiIIScheduleController_5_reset = reset;
  assign MultiIIScheduleController_5_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_5_io_schedules_0 = scheduleDispatch_io_outs_20; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_5_io_schedules_1 = scheduleDispatch_io_outs_21; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_5_io_schedules_2 = scheduleDispatch_io_outs_22; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_5_io_schedules_3 = scheduleDispatch_io_outs_23; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_5_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_6_clock = clock;
  assign MultiIIScheduleController_6_reset = reset;
  assign MultiIIScheduleController_6_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_6_io_schedules_0 = scheduleDispatch_io_outs_24; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_6_io_schedules_1 = scheduleDispatch_io_outs_25; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_6_io_schedules_2 = scheduleDispatch_io_outs_26; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_6_io_schedules_3 = scheduleDispatch_io_outs_27; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_6_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_7_clock = clock;
  assign MultiIIScheduleController_7_reset = reset;
  assign MultiIIScheduleController_7_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_7_io_schedules_0 = scheduleDispatch_io_outs_28; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_7_io_schedules_1 = scheduleDispatch_io_outs_29; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_7_io_schedules_2 = scheduleDispatch_io_outs_30; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_7_io_schedules_3 = scheduleDispatch_io_outs_31; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_7_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_8_clock = clock;
  assign MultiIIScheduleController_8_reset = reset;
  assign MultiIIScheduleController_8_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_8_io_schedules_0 = scheduleDispatch_io_outs_32; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_8_io_schedules_1 = scheduleDispatch_io_outs_33; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_8_io_schedules_2 = scheduleDispatch_io_outs_34; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_8_io_schedules_3 = scheduleDispatch_io_outs_35; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_8_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_9_clock = clock;
  assign MultiIIScheduleController_9_reset = reset;
  assign MultiIIScheduleController_9_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_9_io_schedules_0 = scheduleDispatch_io_outs_36; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_9_io_schedules_1 = scheduleDispatch_io_outs_37; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_9_io_schedules_2 = scheduleDispatch_io_outs_38; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_9_io_schedules_3 = scheduleDispatch_io_outs_39; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_9_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_10_clock = clock;
  assign MultiIIScheduleController_10_reset = reset;
  assign MultiIIScheduleController_10_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_10_io_schedules_0 = scheduleDispatch_io_outs_40; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_10_io_schedules_1 = scheduleDispatch_io_outs_41; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_10_io_schedules_2 = scheduleDispatch_io_outs_42; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_10_io_schedules_3 = scheduleDispatch_io_outs_43; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_10_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_11_clock = clock;
  assign MultiIIScheduleController_11_reset = reset;
  assign MultiIIScheduleController_11_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_11_io_schedules_0 = scheduleDispatch_io_outs_44; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_11_io_schedules_1 = scheduleDispatch_io_outs_45; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_11_io_schedules_2 = scheduleDispatch_io_outs_46; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_11_io_schedules_3 = scheduleDispatch_io_outs_47; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_11_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_12_clock = clock;
  assign MultiIIScheduleController_12_reset = reset;
  assign MultiIIScheduleController_12_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_12_io_schedules_0 = scheduleDispatch_io_outs_48; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_12_io_schedules_1 = scheduleDispatch_io_outs_49; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_12_io_schedules_2 = scheduleDispatch_io_outs_50; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_12_io_schedules_3 = scheduleDispatch_io_outs_51; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_12_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_13_clock = clock;
  assign MultiIIScheduleController_13_reset = reset;
  assign MultiIIScheduleController_13_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_13_io_schedules_0 = scheduleDispatch_io_outs_52; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_13_io_schedules_1 = scheduleDispatch_io_outs_53; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_13_io_schedules_2 = scheduleDispatch_io_outs_54; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_13_io_schedules_3 = scheduleDispatch_io_outs_55; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_13_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_14_clock = clock;
  assign MultiIIScheduleController_14_reset = reset;
  assign MultiIIScheduleController_14_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_14_io_schedules_0 = scheduleDispatch_io_outs_56; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_14_io_schedules_1 = scheduleDispatch_io_outs_57; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_14_io_schedules_2 = scheduleDispatch_io_outs_58; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_14_io_schedules_3 = scheduleDispatch_io_outs_59; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_14_io_II = io_II; // @[TopModule.scala 131:33]
  assign MultiIIScheduleController_15_clock = clock;
  assign MultiIIScheduleController_15_reset = reset;
  assign MultiIIScheduleController_15_io_en = io_en; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_15_io_schedules_0 = scheduleDispatch_io_outs_60; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_15_io_schedules_1 = scheduleDispatch_io_outs_61; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_15_io_schedules_2 = scheduleDispatch_io_outs_62; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_15_io_schedules_3 = scheduleDispatch_io_outs_63; // @[TopModule.scala 133:45]
  assign MultiIIScheduleController_15_io_II = io_II; // @[TopModule.scala 131:33]
  assign RegisterFile_clock = clock;
  assign RegisterFile_reset = reset;
  assign RegisterFile_io_configuration = Dispatch_1_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_io_inputs_0 = Alu_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_1_clock = clock;
  assign RegisterFile_1_reset = reset;
  assign RegisterFile_1_io_configuration = Dispatch_2_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_1_io_inputs_0 = Alu_1_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_2_clock = clock;
  assign RegisterFile_2_reset = reset;
  assign RegisterFile_2_io_configuration = Dispatch_3_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_2_io_inputs_0 = Alu_2_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_3_clock = clock;
  assign RegisterFile_3_reset = reset;
  assign RegisterFile_3_io_configuration = Dispatch_4_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_3_io_inputs_0 = Alu_3_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_4_clock = clock;
  assign RegisterFile_4_reset = reset;
  assign RegisterFile_4_io_configuration = Dispatch_5_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_4_io_inputs_0 = Alu_4_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_5_clock = clock;
  assign RegisterFile_5_reset = reset;
  assign RegisterFile_5_io_configuration = Dispatch_6_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_5_io_inputs_0 = Alu_5_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_6_clock = clock;
  assign RegisterFile_6_reset = reset;
  assign RegisterFile_6_io_configuration = Dispatch_7_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_6_io_inputs_0 = Alu_6_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_7_clock = clock;
  assign RegisterFile_7_reset = reset;
  assign RegisterFile_7_io_configuration = Dispatch_8_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_7_io_inputs_0 = Alu_7_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_8_clock = clock;
  assign RegisterFile_8_reset = reset;
  assign RegisterFile_8_io_configuration = Dispatch_9_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_8_io_inputs_0 = Alu_8_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_9_clock = clock;
  assign RegisterFile_9_reset = reset;
  assign RegisterFile_9_io_configuration = Dispatch_10_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_9_io_inputs_0 = Alu_9_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_10_clock = clock;
  assign RegisterFile_10_reset = reset;
  assign RegisterFile_10_io_configuration = Dispatch_11_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_10_io_inputs_0 = Alu_10_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_11_clock = clock;
  assign RegisterFile_11_reset = reset;
  assign RegisterFile_11_io_configuration = Dispatch_12_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_11_io_inputs_0 = Alu_11_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_12_clock = clock;
  assign RegisterFile_12_reset = reset;
  assign RegisterFile_12_io_configuration = Dispatch_13_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_12_io_inputs_0 = Alu_12_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_13_clock = clock;
  assign RegisterFile_13_reset = reset;
  assign RegisterFile_13_io_configuration = Dispatch_14_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_13_io_inputs_0 = Alu_13_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_14_clock = clock;
  assign RegisterFile_14_reset = reset;
  assign RegisterFile_14_io_configuration = Dispatch_15_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_14_io_inputs_0 = Alu_14_io_outs_0; // @[TopModule.scala 267:60]
  assign RegisterFile_15_clock = clock;
  assign RegisterFile_15_reset = reset;
  assign RegisterFile_15_io_configuration = Dispatch_16_io_outs_1; // @[TopModule.scala 242:22]
  assign RegisterFile_15_io_inputs_0 = Alu_15_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_io_configuration = Dispatch_io_outs_0; // @[TopModule.scala 242:22]
  assign Multiplexer_io_inputs_3 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_io_inputs_2 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_io_inputs_1 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_io_inputs_0 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_1_io_configuration = Dispatch_io_outs_1; // @[TopModule.scala 242:22]
  assign Multiplexer_1_io_inputs_1 = io_inputs_1; // @[TopModule.scala 265:60]
  assign Multiplexer_1_io_inputs_0 = io_inputs_0; // @[TopModule.scala 265:60]
  assign Multiplexer_2_io_configuration = Dispatch_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_2_io_inputs_1 = io_inputs_1; // @[TopModule.scala 265:60]
  assign Multiplexer_2_io_inputs_0 = io_inputs_0; // @[TopModule.scala 265:60]
  assign Multiplexer_3_io_configuration = Dispatch_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_3_io_inputs_1 = io_inputs_1; // @[TopModule.scala 265:60]
  assign Multiplexer_3_io_inputs_0 = io_inputs_0; // @[TopModule.scala 265:60]
  assign Multiplexer_4_io_configuration = Dispatch_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_4_io_inputs_1 = io_inputs_1; // @[TopModule.scala 265:60]
  assign Multiplexer_4_io_inputs_0 = io_inputs_0; // @[TopModule.scala 265:60]
  assign Multiplexer_5_io_configuration = Dispatch_1_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_5_io_inputs_5 = RegisterFile_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_3 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_2 = Multiplexer_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_1 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_5_io_inputs_0 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_6_io_configuration = Dispatch_1_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_6_io_inputs_4 = ConstUnit_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_6_io_inputs_3 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_6_io_inputs_2 = Multiplexer_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_6_io_inputs_1 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_6_io_inputs_0 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_configuration = Dispatch_1_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_7_io_inputs_3 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_2 = Multiplexer_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_1 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_7_io_inputs_0 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_8_io_configuration = Dispatch_1_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_8_io_inputs_1 = Multiplexer_7_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_8_io_inputs_0 = RegisterFile_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_configuration = Dispatch_2_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_9_io_inputs_5 = RegisterFile_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_4 = ConstUnit_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_3 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_2 = Multiplexer_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_1 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_9_io_inputs_0 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_10_io_configuration = Dispatch_2_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_10_io_inputs_4 = ConstUnit_1_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_10_io_inputs_3 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_10_io_inputs_2 = Multiplexer_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_10_io_inputs_1 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_10_io_inputs_0 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_configuration = Dispatch_2_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_11_io_inputs_3 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_2 = Multiplexer_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_1 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_11_io_inputs_0 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_12_io_configuration = Dispatch_2_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_12_io_inputs_1 = Multiplexer_11_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_12_io_inputs_0 = RegisterFile_1_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_configuration = Dispatch_3_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_13_io_inputs_5 = RegisterFile_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_4 = ConstUnit_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_3 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_2 = Multiplexer_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_1 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_13_io_inputs_0 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_14_io_configuration = Dispatch_3_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_14_io_inputs_4 = ConstUnit_2_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_14_io_inputs_3 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_14_io_inputs_2 = Multiplexer_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_14_io_inputs_1 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_14_io_inputs_0 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_configuration = Dispatch_3_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_15_io_inputs_3 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_2 = Multiplexer_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_1 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_15_io_inputs_0 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_16_io_configuration = Dispatch_3_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_16_io_inputs_1 = Multiplexer_15_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_16_io_inputs_0 = RegisterFile_2_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_configuration = Dispatch_4_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_17_io_inputs_5 = RegisterFile_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_4 = ConstUnit_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_3 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_2 = Multiplexer_4_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_1 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_17_io_inputs_0 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_18_io_configuration = Dispatch_4_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_18_io_inputs_4 = ConstUnit_3_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_18_io_inputs_3 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_18_io_inputs_2 = Multiplexer_4_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_18_io_inputs_1 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_18_io_inputs_0 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_19_io_configuration = Dispatch_4_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_19_io_inputs_3 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_19_io_inputs_2 = Multiplexer_4_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_19_io_inputs_1 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_19_io_inputs_0 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_20_io_configuration = Dispatch_4_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_20_io_inputs_1 = Multiplexer_19_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_20_io_inputs_0 = RegisterFile_3_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_21_io_configuration = Dispatch_5_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_21_io_inputs_5 = RegisterFile_4_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_21_io_inputs_4 = ConstUnit_4_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_21_io_inputs_3 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_21_io_inputs_2 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_21_io_inputs_1 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_21_io_inputs_0 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_22_io_configuration = Dispatch_5_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_22_io_inputs_4 = ConstUnit_4_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_22_io_inputs_3 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_22_io_inputs_2 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_22_io_inputs_1 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_22_io_inputs_0 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_23_io_configuration = Dispatch_5_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_23_io_inputs_3 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_23_io_inputs_2 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_23_io_inputs_1 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_23_io_inputs_0 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_24_io_configuration = Dispatch_5_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_24_io_inputs_1 = Multiplexer_23_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_24_io_inputs_0 = RegisterFile_4_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_25_io_configuration = Dispatch_6_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_25_io_inputs_5 = RegisterFile_5_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_25_io_inputs_4 = ConstUnit_5_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_25_io_inputs_3 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_25_io_inputs_2 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_25_io_inputs_1 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_25_io_inputs_0 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_26_io_configuration = Dispatch_6_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_26_io_inputs_4 = ConstUnit_5_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_26_io_inputs_3 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_26_io_inputs_2 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_26_io_inputs_1 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_26_io_inputs_0 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_27_io_configuration = Dispatch_6_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_27_io_inputs_3 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_27_io_inputs_2 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_27_io_inputs_1 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_27_io_inputs_0 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_28_io_configuration = Dispatch_6_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_28_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_28_io_inputs_0 = RegisterFile_5_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_29_io_configuration = Dispatch_7_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_29_io_inputs_5 = RegisterFile_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_29_io_inputs_4 = ConstUnit_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_29_io_inputs_3 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_29_io_inputs_2 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_29_io_inputs_1 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_29_io_inputs_0 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_30_io_configuration = Dispatch_7_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_30_io_inputs_4 = ConstUnit_6_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_30_io_inputs_3 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_30_io_inputs_2 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_30_io_inputs_1 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_30_io_inputs_0 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_31_io_configuration = Dispatch_7_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_31_io_inputs_3 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_31_io_inputs_2 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_31_io_inputs_1 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_31_io_inputs_0 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_32_io_configuration = Dispatch_7_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_32_io_inputs_1 = Multiplexer_31_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_32_io_inputs_0 = RegisterFile_6_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_33_io_configuration = Dispatch_8_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_33_io_inputs_5 = RegisterFile_7_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_33_io_inputs_4 = ConstUnit_7_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_33_io_inputs_3 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_33_io_inputs_2 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_33_io_inputs_1 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_33_io_inputs_0 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_34_io_configuration = Dispatch_8_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_34_io_inputs_4 = ConstUnit_7_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_34_io_inputs_3 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_34_io_inputs_2 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_34_io_inputs_1 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_34_io_inputs_0 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_35_io_configuration = Dispatch_8_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_35_io_inputs_3 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_35_io_inputs_2 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_35_io_inputs_1 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_35_io_inputs_0 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_36_io_configuration = Dispatch_8_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_36_io_inputs_1 = Multiplexer_35_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_36_io_inputs_0 = RegisterFile_7_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_37_io_configuration = Dispatch_9_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_37_io_inputs_5 = RegisterFile_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_37_io_inputs_4 = ConstUnit_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_37_io_inputs_3 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_37_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_37_io_inputs_1 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_37_io_inputs_0 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_38_io_configuration = Dispatch_9_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_38_io_inputs_4 = ConstUnit_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_38_io_inputs_3 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_38_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_38_io_inputs_1 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_38_io_inputs_0 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_39_io_configuration = Dispatch_9_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_39_io_inputs_3 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_39_io_inputs_2 = Multiplexer_24_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_39_io_inputs_1 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_39_io_inputs_0 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_40_io_configuration = Dispatch_9_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_40_io_inputs_1 = Multiplexer_39_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_40_io_inputs_0 = RegisterFile_8_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_41_io_configuration = Dispatch_10_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_41_io_inputs_5 = RegisterFile_9_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_41_io_inputs_4 = ConstUnit_9_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_41_io_inputs_3 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_41_io_inputs_2 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_41_io_inputs_1 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_41_io_inputs_0 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_42_io_configuration = Dispatch_10_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_42_io_inputs_4 = ConstUnit_9_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_42_io_inputs_3 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_42_io_inputs_2 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_42_io_inputs_1 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_42_io_inputs_0 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_43_io_configuration = Dispatch_10_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_43_io_inputs_3 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_43_io_inputs_2 = Multiplexer_28_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_43_io_inputs_1 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_43_io_inputs_0 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_44_io_configuration = Dispatch_10_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_44_io_inputs_1 = Multiplexer_43_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_44_io_inputs_0 = RegisterFile_9_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_45_io_configuration = Dispatch_11_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_45_io_inputs_5 = RegisterFile_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_45_io_inputs_4 = ConstUnit_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_45_io_inputs_3 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_45_io_inputs_2 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_45_io_inputs_1 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_45_io_inputs_0 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_46_io_configuration = Dispatch_11_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_46_io_inputs_4 = ConstUnit_10_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_46_io_inputs_3 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_46_io_inputs_2 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_46_io_inputs_1 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_46_io_inputs_0 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_47_io_configuration = Dispatch_11_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_47_io_inputs_3 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_47_io_inputs_2 = Multiplexer_32_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_47_io_inputs_1 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_47_io_inputs_0 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_48_io_configuration = Dispatch_11_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_48_io_inputs_1 = Multiplexer_47_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_48_io_inputs_0 = RegisterFile_10_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_49_io_configuration = Dispatch_12_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_49_io_inputs_5 = RegisterFile_11_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_49_io_inputs_4 = ConstUnit_11_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_49_io_inputs_3 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_49_io_inputs_2 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_49_io_inputs_1 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_49_io_inputs_0 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_50_io_configuration = Dispatch_12_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_50_io_inputs_4 = ConstUnit_11_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_50_io_inputs_3 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_50_io_inputs_2 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_50_io_inputs_1 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_50_io_inputs_0 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_51_io_configuration = Dispatch_12_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_51_io_inputs_3 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_51_io_inputs_2 = Multiplexer_36_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_51_io_inputs_1 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_51_io_inputs_0 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_52_io_configuration = Dispatch_12_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_52_io_inputs_1 = Multiplexer_51_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_52_io_inputs_0 = RegisterFile_11_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_53_io_configuration = Dispatch_13_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_53_io_inputs_5 = RegisterFile_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_53_io_inputs_4 = ConstUnit_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_53_io_inputs_3 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_53_io_inputs_2 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_53_io_inputs_1 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_53_io_inputs_0 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_54_io_configuration = Dispatch_13_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_54_io_inputs_4 = ConstUnit_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_54_io_inputs_3 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_54_io_inputs_2 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_54_io_inputs_1 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_54_io_inputs_0 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_55_io_configuration = Dispatch_13_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_55_io_inputs_3 = Multiplexer_8_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_55_io_inputs_2 = Multiplexer_40_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_55_io_inputs_1 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_55_io_inputs_0 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_56_io_configuration = Dispatch_13_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_56_io_inputs_1 = Multiplexer_55_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_56_io_inputs_0 = RegisterFile_12_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_57_io_configuration = Dispatch_14_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_57_io_inputs_5 = RegisterFile_13_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_57_io_inputs_4 = ConstUnit_13_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_57_io_inputs_3 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_57_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_57_io_inputs_1 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_57_io_inputs_0 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_58_io_configuration = Dispatch_14_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_58_io_inputs_4 = ConstUnit_13_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_58_io_inputs_3 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_58_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_58_io_inputs_1 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_58_io_inputs_0 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_59_io_configuration = Dispatch_14_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_59_io_inputs_3 = Multiplexer_12_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_59_io_inputs_2 = Multiplexer_44_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_59_io_inputs_1 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_59_io_inputs_0 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_60_io_configuration = Dispatch_14_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_60_io_inputs_1 = Multiplexer_59_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_60_io_inputs_0 = RegisterFile_13_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_61_io_configuration = Dispatch_15_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_61_io_inputs_5 = RegisterFile_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_61_io_inputs_4 = ConstUnit_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_61_io_inputs_3 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_61_io_inputs_2 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_61_io_inputs_1 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_61_io_inputs_0 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_62_io_configuration = Dispatch_15_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_62_io_inputs_4 = ConstUnit_14_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_62_io_inputs_3 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_62_io_inputs_2 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_62_io_inputs_1 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_62_io_inputs_0 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_63_io_configuration = Dispatch_15_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_63_io_inputs_3 = Multiplexer_16_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_63_io_inputs_2 = Multiplexer_48_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_63_io_inputs_1 = Multiplexer_68_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_63_io_inputs_0 = Multiplexer_60_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_64_io_configuration = Dispatch_15_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_64_io_inputs_1 = Multiplexer_63_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_64_io_inputs_0 = RegisterFile_14_io_outs_1; // @[TopModule.scala 267:60]
  assign Multiplexer_65_io_configuration = Dispatch_16_io_outs_2; // @[TopModule.scala 242:22]
  assign Multiplexer_65_io_inputs_5 = RegisterFile_15_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_65_io_inputs_4 = ConstUnit_15_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_65_io_inputs_3 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_65_io_inputs_2 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_65_io_inputs_1 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_65_io_inputs_0 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_66_io_configuration = Dispatch_16_io_outs_3; // @[TopModule.scala 242:22]
  assign Multiplexer_66_io_inputs_4 = ConstUnit_15_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_66_io_inputs_3 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_66_io_inputs_2 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_66_io_inputs_1 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_66_io_inputs_0 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_67_io_configuration = Dispatch_16_io_outs_4; // @[TopModule.scala 242:22]
  assign Multiplexer_67_io_inputs_3 = Multiplexer_20_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_67_io_inputs_2 = Multiplexer_52_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_67_io_inputs_1 = Multiplexer_56_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_67_io_inputs_0 = Multiplexer_64_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_68_io_configuration = Dispatch_16_io_outs_5; // @[TopModule.scala 242:22]
  assign Multiplexer_68_io_inputs_1 = Multiplexer_67_io_outs_0; // @[TopModule.scala 267:60]
  assign Multiplexer_68_io_inputs_0 = RegisterFile_15_io_outs_1; // @[TopModule.scala 267:60]
  assign ConstUnit_io_configuration = Dispatch_1_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_1_io_configuration = Dispatch_2_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_2_io_configuration = Dispatch_3_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_3_io_configuration = Dispatch_4_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_4_io_configuration = Dispatch_5_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_5_io_configuration = Dispatch_6_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_6_io_configuration = Dispatch_7_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_7_io_configuration = Dispatch_8_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_8_io_configuration = Dispatch_9_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_9_io_configuration = Dispatch_10_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_10_io_configuration = Dispatch_11_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_11_io_configuration = Dispatch_12_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_12_io_configuration = Dispatch_13_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_13_io_configuration = Dispatch_14_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_14_io_configuration = Dispatch_15_io_outs_6; // @[TopModule.scala 242:22]
  assign ConstUnit_15_io_configuration = Dispatch_16_io_outs_6; // @[TopModule.scala 242:22]
  assign configControllers_0_clock = clock;
  assign configControllers_0_reset = reset;
  assign configControllers_0_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_0_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_0_io_inConfig = topDispatch_io_outs_0; // @[TopModule.scala 252:38]
  assign Dispatch_io_configuration = configControllers_0_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_1_clock = clock;
  assign configControllers_1_reset = reset;
  assign configControllers_1_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_1_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_1_io_inConfig = topDispatch_io_outs_1; // @[TopModule.scala 252:38]
  assign Dispatch_1_io_configuration = configControllers_1_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_2_clock = clock;
  assign configControllers_2_reset = reset;
  assign configControllers_2_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_2_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_2_io_inConfig = topDispatch_io_outs_2; // @[TopModule.scala 252:38]
  assign Dispatch_2_io_configuration = configControllers_2_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_3_clock = clock;
  assign configControllers_3_reset = reset;
  assign configControllers_3_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_3_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_3_io_inConfig = topDispatch_io_outs_3; // @[TopModule.scala 252:38]
  assign Dispatch_3_io_configuration = configControllers_3_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_4_clock = clock;
  assign configControllers_4_reset = reset;
  assign configControllers_4_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_4_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_4_io_inConfig = topDispatch_io_outs_4; // @[TopModule.scala 252:38]
  assign Dispatch_4_io_configuration = configControllers_4_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_5_clock = clock;
  assign configControllers_5_reset = reset;
  assign configControllers_5_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_5_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_5_io_inConfig = topDispatch_io_outs_5; // @[TopModule.scala 252:38]
  assign Dispatch_5_io_configuration = configControllers_5_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_6_clock = clock;
  assign configControllers_6_reset = reset;
  assign configControllers_6_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_6_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_6_io_inConfig = topDispatch_io_outs_6; // @[TopModule.scala 252:38]
  assign Dispatch_6_io_configuration = configControllers_6_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_7_clock = clock;
  assign configControllers_7_reset = reset;
  assign configControllers_7_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_7_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_7_io_inConfig = topDispatch_io_outs_7; // @[TopModule.scala 252:38]
  assign Dispatch_7_io_configuration = configControllers_7_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_8_clock = clock;
  assign configControllers_8_reset = reset;
  assign configControllers_8_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_8_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_8_io_inConfig = topDispatch_io_outs_8; // @[TopModule.scala 252:38]
  assign Dispatch_8_io_configuration = configControllers_8_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_9_clock = clock;
  assign configControllers_9_reset = reset;
  assign configControllers_9_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_9_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_9_io_inConfig = topDispatch_io_outs_9; // @[TopModule.scala 252:38]
  assign Dispatch_9_io_configuration = configControllers_9_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_10_clock = clock;
  assign configControllers_10_reset = reset;
  assign configControllers_10_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_10_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_10_io_inConfig = topDispatch_io_outs_10; // @[TopModule.scala 252:38]
  assign Dispatch_10_io_configuration = configControllers_10_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_11_clock = clock;
  assign configControllers_11_reset = reset;
  assign configControllers_11_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_11_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_11_io_inConfig = topDispatch_io_outs_11; // @[TopModule.scala 252:38]
  assign Dispatch_11_io_configuration = configControllers_11_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_12_clock = clock;
  assign configControllers_12_reset = reset;
  assign configControllers_12_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_12_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_12_io_inConfig = topDispatch_io_outs_12; // @[TopModule.scala 252:38]
  assign Dispatch_12_io_configuration = configControllers_12_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_13_clock = clock;
  assign configControllers_13_reset = reset;
  assign configControllers_13_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_13_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_13_io_inConfig = topDispatch_io_outs_13; // @[TopModule.scala 252:38]
  assign Dispatch_13_io_configuration = configControllers_13_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_14_clock = clock;
  assign configControllers_14_reset = reset;
  assign configControllers_14_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_14_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_14_io_inConfig = topDispatch_io_outs_14; // @[TopModule.scala 252:38]
  assign Dispatch_14_io_configuration = configControllers_14_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_15_clock = clock;
  assign configControllers_15_reset = reset;
  assign configControllers_15_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_15_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_15_io_inConfig = topDispatch_io_outs_15; // @[TopModule.scala 252:38]
  assign Dispatch_15_io_configuration = configControllers_15_io_outConfig; // @[TopModule.scala 245:31]
  assign configControllers_16_clock = clock;
  assign configControllers_16_reset = reset;
  assign configControllers_16_io_en = io_enConfig; // @[TopModule.scala 236:28]
  assign configControllers_16_io_II = io_II; // @[TopModule.scala 235:28]
  assign configControllers_16_io_inConfig = topDispatch_io_outs_16; // @[TopModule.scala 252:38]
  assign Dispatch_16_io_configuration = configControllers_16_io_outConfig; // @[TopModule.scala 245:31]
  assign topDispatch_io_configuration = io_configuration; // @[TopModule.scala 250:32]
endmodule
