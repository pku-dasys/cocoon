module Dispatch(
  input        io_en,
  output [8:0] io_outs_144
);
  assign io_outs_144 = io_en ? 9'h10 : 9'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module RegNextN(
  input         clock,
  input         reset,
  input  [3:0]  io_latency,
  input  [31:0] io_input,
  output [31:0] io_out
);
  reg [31:0] regArray_0; // @[BasicChiselModules.scala 18:25]
  reg [31:0] _RAND_0;
  reg [31:0] regArray_1; // @[BasicChiselModules.scala 18:25]
  reg [31:0] _RAND_1;
  reg [31:0] regArray_2; // @[BasicChiselModules.scala 18:25]
  reg [31:0] _RAND_2;
  wire  _T_1; // @[BasicChiselModules.scala 23:19]
  wire [3:0] _T_3; // @[BasicChiselModules.scala 24:35]
  wire [1:0] _T_4;
  wire [31:0] _GEN_1; // @[BasicChiselModules.scala 24:12]
  wire [31:0] _GEN_2; // @[BasicChiselModules.scala 24:12]
  assign _T_1 = io_latency > 4'h0; // @[BasicChiselModules.scala 23:19]
  assign _T_3 = io_latency - 4'h1; // @[BasicChiselModules.scala 24:35]
  assign _T_4 = _T_3[1:0];
  assign _GEN_1 = 2'h1 == _T_4 ? regArray_1 : regArray_0; // @[BasicChiselModules.scala 24:12]
  assign _GEN_2 = 2'h2 == _T_4 ? regArray_2 : _GEN_1; // @[BasicChiselModules.scala 24:12]
  assign io_out = _T_1 ? _GEN_2 : io_input; // @[BasicChiselModules.scala 24:12 BasicChiselModules.scala 26:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regArray_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regArray_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regArray_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regArray_0 <= 32'h0;
    end else begin
      regArray_0 <= io_input;
    end
    if (reset) begin
      regArray_1 <= 32'h0;
    end else begin
      regArray_1 <= regArray_0;
    end
    if (reset) begin
      regArray_2 <= 32'h0;
    end else begin
      regArray_2 <= regArray_1;
    end
  end
endmodule
module SyncScheduleController(
  input         clock,
  input         reset,
  input  [4:0]  io_skewing,
  input  [31:0] io_input0,
  input  [31:0] io_input1,
  output [31:0] io_skewedInput0,
  output [31:0] io_skewedInput1
);
  wire  regNextN_clock; // @[BasicChiselModules.scala 39:24]
  wire  regNextN_reset; // @[BasicChiselModules.scala 39:24]
  wire [3:0] regNextN_io_latency; // @[BasicChiselModules.scala 39:24]
  wire [31:0] regNextN_io_input; // @[BasicChiselModules.scala 39:24]
  wire [31:0] regNextN_io_out; // @[BasicChiselModules.scala 39:24]
  wire  signal; // @[BasicChiselModules.scala 41:26]
  RegNextN regNextN ( // @[BasicChiselModules.scala 39:24]
    .clock(regNextN_clock),
    .reset(regNextN_reset),
    .io_latency(regNextN_io_latency),
    .io_input(regNextN_io_input),
    .io_out(regNextN_io_out)
  );
  assign signal = io_skewing[4]; // @[BasicChiselModules.scala 41:26]
  assign io_skewedInput0 = signal ? regNextN_io_out : io_input0; // @[BasicChiselModules.scala 46:21 BasicChiselModules.scala 51:21]
  assign io_skewedInput1 = signal ? io_input1 : regNextN_io_out; // @[BasicChiselModules.scala 47:21 BasicChiselModules.scala 50:21]
  assign regNextN_clock = clock;
  assign regNextN_reset = reset;
  assign regNextN_io_latency = io_skewing[3:0]; // @[BasicChiselModules.scala 42:23]
  assign regNextN_io_input = signal ? io_input0 : io_input1; // @[BasicChiselModules.scala 45:23 BasicChiselModules.scala 49:23]
endmodule
module Alu(
  input         clock,
  input         reset,
  input         io_en,
  input  [4:0]  io_skewing,
  input  [3:0]  io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  syncScheduleController_clock; // @[BasicChiselModules.scala 198:38]
  wire  syncScheduleController_reset; // @[BasicChiselModules.scala 198:38]
  wire [4:0] syncScheduleController_io_skewing; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_input0; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_input1; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_skewedInput0; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 198:38]
  wire [5:0] shamt; // @[BasicChiselModules.scala 207:22]
  wire [31:0] _T_1; // @[BasicChiselModules.scala 176:55]
  wire [31:0] _T_3; // @[BasicChiselModules.scala 177:55]
  wire [31:0] _T_4; // @[BasicChiselModules.scala 178:55]
  wire [31:0] _T_5; // @[BasicChiselModules.scala 179:54]
  wire [31:0] _T_6; // @[BasicChiselModules.scala 180:55]
  wire [63:0] _T_7; // @[BasicChiselModules.scala 181:55]
  wire [94:0] _GEN_1; // @[BasicChiselModules.scala 183:56]
  wire [94:0] _T_8; // @[BasicChiselModules.scala 183:56]
  wire [31:0] _T_9; // @[BasicChiselModules.scala 186:56]
  wire [31:0] _T_10; // @[BasicChiselModules.scala 188:57]
  wire [31:0] _T_11; // @[BasicChiselModules.scala 188:64]
  wire [31:0] _T_12; // @[BasicChiselModules.scala 188:74]
  wire [31:0] _T_13; // @[BasicChiselModules.scala 189:55]
  wire [31:0] _T_15; // @[Mux.scala 68:16]
  wire  _T_16; // @[Mux.scala 68:19]
  wire [31:0] _T_17; // @[Mux.scala 68:16]
  wire  _T_18; // @[Mux.scala 68:19]
  wire [31:0] _T_19; // @[Mux.scala 68:16]
  wire  _T_20; // @[Mux.scala 68:19]
  wire [31:0] _T_21; // @[Mux.scala 68:16]
  wire  _T_22; // @[Mux.scala 68:19]
  wire [31:0] _T_23; // @[Mux.scala 68:16]
  wire  _T_24; // @[Mux.scala 68:19]
  wire [94:0] _T_25; // @[Mux.scala 68:16]
  wire  _T_26; // @[Mux.scala 68:19]
  wire [94:0] _T_27; // @[Mux.scala 68:16]
  wire  _T_28; // @[Mux.scala 68:19]
  wire [94:0] _T_29; // @[Mux.scala 68:16]
  wire  _T_30; // @[Mux.scala 68:19]
  wire [94:0] _T_31; // @[Mux.scala 68:16]
  wire  _T_32; // @[Mux.scala 68:19]
  wire [94:0] _T_33; // @[Mux.scala 68:16]
  wire  _T_34; // @[Mux.scala 68:19]
  wire [94:0] _T_35; // @[Mux.scala 68:16]
  wire  _T_36; // @[Mux.scala 68:19]
  wire [94:0] _T_37; // @[Mux.scala 68:16]
  wire [94:0] _GEN_0; // @[BasicChiselModules.scala 211:14]
  SyncScheduleController syncScheduleController ( // @[BasicChiselModules.scala 198:38]
    .clock(syncScheduleController_clock),
    .reset(syncScheduleController_reset),
    .io_skewing(syncScheduleController_io_skewing),
    .io_input0(syncScheduleController_io_input0),
    .io_input1(syncScheduleController_io_input1),
    .io_skewedInput0(syncScheduleController_io_skewedInput0),
    .io_skewedInput1(syncScheduleController_io_skewedInput1)
  );
  assign shamt = syncScheduleController_io_skewedInput1[5:0]; // @[BasicChiselModules.scala 207:22]
  assign _T_1 = syncScheduleController_io_skewedInput0 + syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 176:55]
  assign _T_3 = syncScheduleController_io_skewedInput0 - syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 177:55]
  assign _T_4 = syncScheduleController_io_skewedInput0 & syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 178:55]
  assign _T_5 = syncScheduleController_io_skewedInput0 | syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 179:54]
  assign _T_6 = syncScheduleController_io_skewedInput0 ^ syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 180:55]
  assign _T_7 = syncScheduleController_io_skewedInput0 * syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 181:55]
  assign _GEN_1 = {{63'd0}, syncScheduleController_io_skewedInput0}; // @[BasicChiselModules.scala 183:56]
  assign _T_8 = _GEN_1 << shamt; // @[BasicChiselModules.scala 183:56]
  assign _T_9 = syncScheduleController_io_skewedInput0 >> shamt; // @[BasicChiselModules.scala 186:56]
  assign _T_10 = $signed(syncScheduleController_io_skewedInput0); // @[BasicChiselModules.scala 188:57]
  assign _T_11 = $signed(_T_10) >>> shamt; // @[BasicChiselModules.scala 188:64]
  assign _T_12 = $unsigned(_T_11); // @[BasicChiselModules.scala 188:74]
  assign _T_13 = syncScheduleController_io_skewedInput0 / syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 189:55]
  assign _T_15 = syncScheduleController_io_skewedInput1; // @[Mux.scala 68:16]
  assign _T_16 = 4'hc == io_configuration; // @[Mux.scala 68:19]
  assign _T_17 = _T_16 ? syncScheduleController_io_skewedInput0 : _T_15; // @[Mux.scala 68:16]
  assign _T_18 = 4'hb == io_configuration; // @[Mux.scala 68:19]
  assign _T_19 = _T_18 ? _T_13 : _T_17; // @[Mux.scala 68:16]
  assign _T_20 = 4'ha == io_configuration; // @[Mux.scala 68:19]
  assign _T_21 = _T_20 ? _T_12 : _T_19; // @[Mux.scala 68:16]
  assign _T_22 = 4'h9 == io_configuration; // @[Mux.scala 68:19]
  assign _T_23 = _T_22 ? _T_9 : _T_21; // @[Mux.scala 68:16]
  assign _T_24 = 4'h7 == io_configuration; // @[Mux.scala 68:19]
  assign _T_25 = _T_24 ? _T_8 : {{63'd0}, _T_23}; // @[Mux.scala 68:16]
  assign _T_26 = 4'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_27 = _T_26 ? {{31'd0}, _T_7} : _T_25; // @[Mux.scala 68:16]
  assign _T_28 = 4'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_29 = _T_28 ? {{63'd0}, _T_6} : _T_27; // @[Mux.scala 68:16]
  assign _T_30 = 4'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_31 = _T_30 ? {{63'd0}, _T_5} : _T_29; // @[Mux.scala 68:16]
  assign _T_32 = 4'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_33 = _T_32 ? {{63'd0}, _T_4} : _T_31; // @[Mux.scala 68:16]
  assign _T_34 = 4'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_35 = _T_34 ? {{63'd0}, _T_3} : _T_33; // @[Mux.scala 68:16]
  assign _T_36 = 4'h0 == io_configuration; // @[Mux.scala 68:19]
  assign _T_37 = _T_36 ? {{63'd0}, _T_1} : _T_35; // @[Mux.scala 68:16]
  assign _GEN_0 = io_en ? _T_37 : 95'h0; // @[BasicChiselModules.scala 211:14]
  assign io_outs_0 = _GEN_0[31:0]; // @[BasicChiselModules.scala 212:9 BasicChiselModules.scala 229:11]
  assign syncScheduleController_clock = clock;
  assign syncScheduleController_reset = reset;
  assign syncScheduleController_io_skewing = io_skewing; // @[BasicChiselModules.scala 202:37]
  assign syncScheduleController_io_input0 = io_inputs_0; // @[BasicChiselModules.scala 199:36]
  assign syncScheduleController_io_input1 = io_inputs_1; // @[BasicChiselModules.scala 200:36]
endmodule
module Alu_4(
  input         clock,
  input         reset,
  input         io_en,
  input  [4:0]  io_skewing,
  input  [3:0]  io_configuration,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  syncScheduleController_clock; // @[BasicChiselModules.scala 198:38]
  wire  syncScheduleController_reset; // @[BasicChiselModules.scala 198:38]
  wire [4:0] syncScheduleController_io_skewing; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_input0; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_input1; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_skewedInput0; // @[BasicChiselModules.scala 198:38]
  wire [31:0] syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 198:38]
  wire [31:0] _T_1; // @[BasicChiselModules.scala 176:55]
  wire [63:0] _T_2; // @[BasicChiselModules.scala 181:55]
  wire [31:0] _T_4; // @[Mux.scala 68:16]
  wire  _T_5; // @[Mux.scala 68:19]
  wire [31:0] _T_6; // @[Mux.scala 68:16]
  wire  _T_7; // @[Mux.scala 68:19]
  wire [63:0] _T_8; // @[Mux.scala 68:16]
  wire  _T_9; // @[Mux.scala 68:19]
  wire [63:0] _T_10; // @[Mux.scala 68:16]
  wire [63:0] _GEN_0; // @[BasicChiselModules.scala 211:14]
  SyncScheduleController syncScheduleController ( // @[BasicChiselModules.scala 198:38]
    .clock(syncScheduleController_clock),
    .reset(syncScheduleController_reset),
    .io_skewing(syncScheduleController_io_skewing),
    .io_input0(syncScheduleController_io_input0),
    .io_input1(syncScheduleController_io_input1),
    .io_skewedInput0(syncScheduleController_io_skewedInput0),
    .io_skewedInput1(syncScheduleController_io_skewedInput1)
  );
  assign _T_1 = syncScheduleController_io_skewedInput0 + syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 176:55]
  assign _T_2 = syncScheduleController_io_skewedInput0 * syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 181:55]
  assign _T_4 = syncScheduleController_io_skewedInput1; // @[Mux.scala 68:16]
  assign _T_5 = 4'hc == io_configuration; // @[Mux.scala 68:19]
  assign _T_6 = _T_5 ? syncScheduleController_io_skewedInput0 : _T_4; // @[Mux.scala 68:16]
  assign _T_7 = 4'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_8 = _T_7 ? _T_2 : {{32'd0}, _T_6}; // @[Mux.scala 68:16]
  assign _T_9 = 4'h0 == io_configuration; // @[Mux.scala 68:19]
  assign _T_10 = _T_9 ? {{32'd0}, _T_1} : _T_8; // @[Mux.scala 68:16]
  assign _GEN_0 = io_en ? _T_10 : 64'h0; // @[BasicChiselModules.scala 211:14]
  assign io_outs_0 = _GEN_0[31:0]; // @[BasicChiselModules.scala 212:9 BasicChiselModules.scala 229:11]
  assign syncScheduleController_clock = clock;
  assign syncScheduleController_reset = reset;
  assign syncScheduleController_io_skewing = io_skewing; // @[BasicChiselModules.scala 202:37]
  assign syncScheduleController_io_input0 = io_inputs_0; // @[BasicChiselModules.scala 199:36]
  assign syncScheduleController_io_input1 = io_inputs_1; // @[BasicChiselModules.scala 200:36]
endmodule
module ScheduleController(
  input        clock,
  input        reset,
  input        io_en,
  input  [3:0] io_waitCycle,
  output       io_valid
);
  reg  state; // @[BasicChiselModules.scala 107:22]
  reg [31:0] _RAND_0;
  reg [3:0] cycleReg; // @[BasicChiselModules.scala 108:21]
  reg [31:0] _RAND_1;
  wire  _T; // @[BasicChiselModules.scala 110:25]
  wire  _T_2; // @[BasicChiselModules.scala 113:16]
  wire [3:0] _T_5; // @[BasicChiselModules.scala 117:30]
  wire  _GEN_0; // @[BasicChiselModules.scala 114:38]
  wire  _GEN_2; // @[BasicChiselModules.scala 113:27]
  wire  _GEN_4; // @[BasicChiselModules.scala 112:14]
  assign _T = cycleReg == io_waitCycle; // @[BasicChiselModules.scala 110:25]
  assign _T_2 = state == 1'h0; // @[BasicChiselModules.scala 113:16]
  assign _T_5 = cycleReg + 4'h1; // @[BasicChiselModules.scala 117:30]
  assign _GEN_0 = _T | state; // @[BasicChiselModules.scala 114:38]
  assign _GEN_2 = _T_2 ? _GEN_0 : state; // @[BasicChiselModules.scala 113:27]
  assign _GEN_4 = io_en & _GEN_2; // @[BasicChiselModules.scala 112:14]
  assign io_valid = _T & io_en; // @[BasicChiselModules.scala 110:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_4;
    end
    if (io_en) begin
      if (_T_2) begin
        if (!(_T)) begin
          cycleReg <= _T_5;
        end
      end
    end else begin
      cycleReg <= 4'h0;
    end
  end
endmodule
module MultiIIScheduleController(
  input        clock,
  input        reset,
  input        io_en,
  input  [8:0] io_schedules_0,
  input  [2:0] io_II,
  output       io_valid,
  output [4:0] io_skewing
);
  wire  ScheduleController_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_io_valid; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_1_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_1_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_1_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_1_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_1_io_valid; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_2_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_2_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_2_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_2_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_2_io_valid; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_3_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_3_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_3_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_3_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_3_io_valid; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_4_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_4_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_4_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_4_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_4_io_valid; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_5_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_5_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_5_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_5_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_5_io_valid; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_6_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_6_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_6_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_6_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_6_io_valid; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_7_clock; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_7_reset; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_7_io_en; // @[BasicChiselModules.scala 134:77]
  wire [3:0] ScheduleController_7_io_waitCycle; // @[BasicChiselModules.scala 134:77]
  wire  ScheduleController_7_io_valid; // @[BasicChiselModules.scala 134:77]
  reg  validRegs_0; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_0;
  reg  validRegs_1; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_1;
  reg  validRegs_2; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_2;
  reg  validRegs_3; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_3;
  reg  validRegs_4; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_4;
  reg  validRegs_5; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_5;
  reg  validRegs_6; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_6;
  reg  validRegs_7; // @[BasicChiselModules.scala 135:26]
  reg [31:0] _RAND_7;
  reg [2:0] cycleReg; // @[BasicChiselModules.scala 136:25]
  reg [31:0] _RAND_8;
  wire  _GEN_1; // @[BasicChiselModules.scala 145:12]
  wire  _GEN_2; // @[BasicChiselModules.scala 145:12]
  wire  _GEN_3; // @[BasicChiselModules.scala 145:12]
  wire  _GEN_4; // @[BasicChiselModules.scala 145:12]
  wire  _GEN_5; // @[BasicChiselModules.scala 145:12]
  wire  _GEN_6; // @[BasicChiselModules.scala 145:12]
  wire [8:0] _GEN_9; // @[BasicChiselModules.scala 146:39]
  wire [8:0] _GEN_10; // @[BasicChiselModules.scala 146:39]
  wire [8:0] _GEN_11; // @[BasicChiselModules.scala 146:39]
  wire [8:0] _GEN_12; // @[BasicChiselModules.scala 146:39]
  wire [8:0] _GEN_13; // @[BasicChiselModules.scala 146:39]
  wire [8:0] _GEN_14; // @[BasicChiselModules.scala 146:39]
  wire [8:0] _GEN_15; // @[BasicChiselModules.scala 146:39]
  wire [2:0] _T_12; // @[BasicChiselModules.scala 149:29]
  wire  _T_13; // @[BasicChiselModules.scala 149:19]
  wire [2:0] _T_15; // @[BasicChiselModules.scala 152:28]
  ScheduleController ScheduleController ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_clock),
    .reset(ScheduleController_reset),
    .io_en(ScheduleController_io_en),
    .io_waitCycle(ScheduleController_io_waitCycle),
    .io_valid(ScheduleController_io_valid)
  );
  ScheduleController ScheduleController_1 ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_1_clock),
    .reset(ScheduleController_1_reset),
    .io_en(ScheduleController_1_io_en),
    .io_waitCycle(ScheduleController_1_io_waitCycle),
    .io_valid(ScheduleController_1_io_valid)
  );
  ScheduleController ScheduleController_2 ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_2_clock),
    .reset(ScheduleController_2_reset),
    .io_en(ScheduleController_2_io_en),
    .io_waitCycle(ScheduleController_2_io_waitCycle),
    .io_valid(ScheduleController_2_io_valid)
  );
  ScheduleController ScheduleController_3 ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_3_clock),
    .reset(ScheduleController_3_reset),
    .io_en(ScheduleController_3_io_en),
    .io_waitCycle(ScheduleController_3_io_waitCycle),
    .io_valid(ScheduleController_3_io_valid)
  );
  ScheduleController ScheduleController_4 ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_4_clock),
    .reset(ScheduleController_4_reset),
    .io_en(ScheduleController_4_io_en),
    .io_waitCycle(ScheduleController_4_io_waitCycle),
    .io_valid(ScheduleController_4_io_valid)
  );
  ScheduleController ScheduleController_5 ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_5_clock),
    .reset(ScheduleController_5_reset),
    .io_en(ScheduleController_5_io_en),
    .io_waitCycle(ScheduleController_5_io_waitCycle),
    .io_valid(ScheduleController_5_io_valid)
  );
  ScheduleController ScheduleController_6 ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_6_clock),
    .reset(ScheduleController_6_reset),
    .io_en(ScheduleController_6_io_en),
    .io_waitCycle(ScheduleController_6_io_waitCycle),
    .io_valid(ScheduleController_6_io_valid)
  );
  ScheduleController ScheduleController_7 ( // @[BasicChiselModules.scala 134:77]
    .clock(ScheduleController_7_clock),
    .reset(ScheduleController_7_reset),
    .io_en(ScheduleController_7_io_en),
    .io_waitCycle(ScheduleController_7_io_waitCycle),
    .io_valid(ScheduleController_7_io_valid)
  );
  assign _GEN_1 = 3'h1 == cycleReg ? validRegs_1 : validRegs_0; // @[BasicChiselModules.scala 145:12]
  assign _GEN_2 = 3'h2 == cycleReg ? validRegs_2 : _GEN_1; // @[BasicChiselModules.scala 145:12]
  assign _GEN_3 = 3'h3 == cycleReg ? validRegs_3 : _GEN_2; // @[BasicChiselModules.scala 145:12]
  assign _GEN_4 = 3'h4 == cycleReg ? validRegs_4 : _GEN_3; // @[BasicChiselModules.scala 145:12]
  assign _GEN_5 = 3'h5 == cycleReg ? validRegs_5 : _GEN_4; // @[BasicChiselModules.scala 145:12]
  assign _GEN_6 = 3'h6 == cycleReg ? validRegs_6 : _GEN_5; // @[BasicChiselModules.scala 145:12]
  assign _GEN_9 = 3'h1 == cycleReg ? 9'h0 : io_schedules_0; // @[BasicChiselModules.scala 146:39]
  assign _GEN_10 = 3'h2 == cycleReg ? 9'h0 : _GEN_9; // @[BasicChiselModules.scala 146:39]
  assign _GEN_11 = 3'h3 == cycleReg ? 9'h0 : _GEN_10; // @[BasicChiselModules.scala 146:39]
  assign _GEN_12 = 3'h4 == cycleReg ? 9'h0 : _GEN_11; // @[BasicChiselModules.scala 146:39]
  assign _GEN_13 = 3'h5 == cycleReg ? 9'h0 : _GEN_12; // @[BasicChiselModules.scala 146:39]
  assign _GEN_14 = 3'h6 == cycleReg ? 9'h0 : _GEN_13; // @[BasicChiselModules.scala 146:39]
  assign _GEN_15 = 3'h7 == cycleReg ? 9'h0 : _GEN_14; // @[BasicChiselModules.scala 146:39]
  assign _T_12 = io_II - 3'h1; // @[BasicChiselModules.scala 149:29]
  assign _T_13 = cycleReg == _T_12; // @[BasicChiselModules.scala 149:19]
  assign _T_15 = cycleReg + 3'h1; // @[BasicChiselModules.scala 152:28]
  assign io_valid = 3'h7 == cycleReg ? validRegs_7 : _GEN_6; // @[BasicChiselModules.scala 145:12]
  assign io_skewing = _GEN_15[8:4]; // @[BasicChiselModules.scala 146:14]
  assign ScheduleController_clock = clock;
  assign ScheduleController_reset = reset;
  assign ScheduleController_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_io_waitCycle = io_schedules_0[3:0]; // @[BasicChiselModules.scala 141:37]
  assign ScheduleController_1_clock = clock;
  assign ScheduleController_1_reset = reset;
  assign ScheduleController_1_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_1_io_waitCycle = 4'h0; // @[BasicChiselModules.scala 141:37]
  assign ScheduleController_2_clock = clock;
  assign ScheduleController_2_reset = reset;
  assign ScheduleController_2_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_2_io_waitCycle = 4'h0; // @[BasicChiselModules.scala 141:37]
  assign ScheduleController_3_clock = clock;
  assign ScheduleController_3_reset = reset;
  assign ScheduleController_3_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_3_io_waitCycle = 4'h0; // @[BasicChiselModules.scala 141:37]
  assign ScheduleController_4_clock = clock;
  assign ScheduleController_4_reset = reset;
  assign ScheduleController_4_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_4_io_waitCycle = 4'h0; // @[BasicChiselModules.scala 141:37]
  assign ScheduleController_5_clock = clock;
  assign ScheduleController_5_reset = reset;
  assign ScheduleController_5_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_5_io_waitCycle = 4'h0; // @[BasicChiselModules.scala 141:37]
  assign ScheduleController_6_clock = clock;
  assign ScheduleController_6_reset = reset;
  assign ScheduleController_6_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_6_io_waitCycle = 4'h0; // @[BasicChiselModules.scala 141:37]
  assign ScheduleController_7_clock = clock;
  assign ScheduleController_7_reset = reset;
  assign ScheduleController_7_io_en = io_en; // @[BasicChiselModules.scala 140:30]
  assign ScheduleController_7_io_waitCycle = 4'h0; // @[BasicChiselModules.scala 141:37]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validRegs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  validRegs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  validRegs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  validRegs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  validRegs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  validRegs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  validRegs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  validRegs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  cycleReg = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      validRegs_0 <= 1'h0;
    end else begin
      validRegs_0 <= ScheduleController_io_valid;
    end
    if (reset) begin
      validRegs_1 <= 1'h0;
    end else begin
      validRegs_1 <= ScheduleController_1_io_valid;
    end
    if (reset) begin
      validRegs_2 <= 1'h0;
    end else begin
      validRegs_2 <= ScheduleController_2_io_valid;
    end
    if (reset) begin
      validRegs_3 <= 1'h0;
    end else begin
      validRegs_3 <= ScheduleController_3_io_valid;
    end
    if (reset) begin
      validRegs_4 <= 1'h0;
    end else begin
      validRegs_4 <= ScheduleController_4_io_valid;
    end
    if (reset) begin
      validRegs_5 <= 1'h0;
    end else begin
      validRegs_5 <= ScheduleController_5_io_valid;
    end
    if (reset) begin
      validRegs_6 <= 1'h0;
    end else begin
      validRegs_6 <= ScheduleController_6_io_valid;
    end
    if (reset) begin
      validRegs_7 <= 1'h0;
    end else begin
      validRegs_7 <= ScheduleController_7_io_valid;
    end
    if (reset) begin
      cycleReg <= 3'h7;
    end else if (io_en) begin
      if (_T_13) begin
        cycleReg <= 3'h0;
      end else begin
        cycleReg <= _T_15;
      end
    end
  end
endmodule
module Dispatch_1(
  input         io_en,
  input  [35:0] io_configuration,
  output [2:0]  io_outs_11,
  output [2:0]  io_outs_10,
  output [2:0]  io_outs_9,
  output [2:0]  io_outs_8,
  output [2:0]  io_outs_7,
  output [2:0]  io_outs_6,
  output [2:0]  io_outs_5,
  output [2:0]  io_outs_4,
  output [2:0]  io_outs_3,
  output [2:0]  io_outs_2,
  output [2:0]  io_outs_1,
  output [2:0]  io_outs_0
);
  wire [2:0] _T; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_1; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_2; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_3; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_4; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_5; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_6; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_7; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_8; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_9; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_10; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_11; // @[BasicChiselModules.scala 409:37]
  assign _T = io_configuration[2:0]; // @[BasicChiselModules.scala 409:37]
  assign _T_1 = io_configuration[5:3]; // @[BasicChiselModules.scala 409:37]
  assign _T_2 = io_configuration[8:6]; // @[BasicChiselModules.scala 409:37]
  assign _T_3 = io_configuration[11:9]; // @[BasicChiselModules.scala 409:37]
  assign _T_4 = io_configuration[14:12]; // @[BasicChiselModules.scala 409:37]
  assign _T_5 = io_configuration[17:15]; // @[BasicChiselModules.scala 409:37]
  assign _T_6 = io_configuration[20:18]; // @[BasicChiselModules.scala 409:37]
  assign _T_7 = io_configuration[23:21]; // @[BasicChiselModules.scala 409:37]
  assign _T_8 = io_configuration[26:24]; // @[BasicChiselModules.scala 409:37]
  assign _T_9 = io_configuration[29:27]; // @[BasicChiselModules.scala 409:37]
  assign _T_10 = io_configuration[32:30]; // @[BasicChiselModules.scala 409:37]
  assign _T_11 = io_configuration[35:33]; // @[BasicChiselModules.scala 409:37]
  assign io_outs_11 = io_en ? _T_11 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_10 = io_en ? _T_10 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_9 = io_en ? _T_9 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_8 = io_en ? _T_8 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_7 = io_en ? _T_7 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_6 = io_en ? _T_6 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_5 = io_en ? _T_5 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_4 = io_en ? _T_4 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_3 = io_en ? _T_3 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_2 = io_en ? _T_2 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_1 = io_en ? _T_1 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_0 = io_en ? _T : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module RegisterFiles(
  input         clock,
  input         reset,
  input         io_en,
  input  [35:0] io_configuration,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_7,
  output [31:0] io_outs_6,
  output [31:0] io_outs_5,
  output [31:0] io_outs_4,
  output [31:0] io_outs_3,
  output [31:0] io_outs_2,
  output [31:0] io_outs_1,
  output [31:0] io_outs_0
);
  wire  dispatch_io_en; // @[BasicChiselModules.scala 275:24]
  wire [35:0] dispatch_io_configuration; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_11; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_10; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_9; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_8; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_7; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_6; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_5; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_4; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_3; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_2; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_1; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_outs_0; // @[BasicChiselModules.scala 275:24]
  reg [31:0] regs_0; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_7;
  wire [31:0] _GEN_33; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_34; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_35; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_36; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_37; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_38; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_39; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_41; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_42; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_43; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_44; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_45; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_46; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_47; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_49; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_50; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_51; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_52; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_53; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_54; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_55; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_57; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_58; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_59; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_60; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_61; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_62; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_63; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_65; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_66; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_67; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_68; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_69; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_70; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_71; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_73; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_74; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_75; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_76; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_77; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_78; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_79; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_81; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_82; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_83; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_84; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_85; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_86; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_87; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_89; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_90; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_91; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_92; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_93; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_94; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_95; // @[BasicChiselModules.scala 292:18]
  Dispatch_1 dispatch ( // @[BasicChiselModules.scala 275:24]
    .io_en(dispatch_io_en),
    .io_configuration(dispatch_io_configuration),
    .io_outs_11(dispatch_io_outs_11),
    .io_outs_10(dispatch_io_outs_10),
    .io_outs_9(dispatch_io_outs_9),
    .io_outs_8(dispatch_io_outs_8),
    .io_outs_7(dispatch_io_outs_7),
    .io_outs_6(dispatch_io_outs_6),
    .io_outs_5(dispatch_io_outs_5),
    .io_outs_4(dispatch_io_outs_4),
    .io_outs_3(dispatch_io_outs_3),
    .io_outs_2(dispatch_io_outs_2),
    .io_outs_1(dispatch_io_outs_1),
    .io_outs_0(dispatch_io_outs_0)
  );
  assign _GEN_33 = 3'h1 == dispatch_io_outs_4 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_34 = 3'h2 == dispatch_io_outs_4 ? regs_2 : _GEN_33; // @[BasicChiselModules.scala 292:18]
  assign _GEN_35 = 3'h3 == dispatch_io_outs_4 ? regs_3 : _GEN_34; // @[BasicChiselModules.scala 292:18]
  assign _GEN_36 = 3'h4 == dispatch_io_outs_4 ? regs_4 : _GEN_35; // @[BasicChiselModules.scala 292:18]
  assign _GEN_37 = 3'h5 == dispatch_io_outs_4 ? regs_5 : _GEN_36; // @[BasicChiselModules.scala 292:18]
  assign _GEN_38 = 3'h6 == dispatch_io_outs_4 ? regs_6 : _GEN_37; // @[BasicChiselModules.scala 292:18]
  assign _GEN_39 = 3'h7 == dispatch_io_outs_4 ? regs_7 : _GEN_38; // @[BasicChiselModules.scala 292:18]
  assign _GEN_41 = 3'h1 == dispatch_io_outs_5 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_42 = 3'h2 == dispatch_io_outs_5 ? regs_2 : _GEN_41; // @[BasicChiselModules.scala 292:18]
  assign _GEN_43 = 3'h3 == dispatch_io_outs_5 ? regs_3 : _GEN_42; // @[BasicChiselModules.scala 292:18]
  assign _GEN_44 = 3'h4 == dispatch_io_outs_5 ? regs_4 : _GEN_43; // @[BasicChiselModules.scala 292:18]
  assign _GEN_45 = 3'h5 == dispatch_io_outs_5 ? regs_5 : _GEN_44; // @[BasicChiselModules.scala 292:18]
  assign _GEN_46 = 3'h6 == dispatch_io_outs_5 ? regs_6 : _GEN_45; // @[BasicChiselModules.scala 292:18]
  assign _GEN_47 = 3'h7 == dispatch_io_outs_5 ? regs_7 : _GEN_46; // @[BasicChiselModules.scala 292:18]
  assign _GEN_49 = 3'h1 == dispatch_io_outs_6 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_50 = 3'h2 == dispatch_io_outs_6 ? regs_2 : _GEN_49; // @[BasicChiselModules.scala 292:18]
  assign _GEN_51 = 3'h3 == dispatch_io_outs_6 ? regs_3 : _GEN_50; // @[BasicChiselModules.scala 292:18]
  assign _GEN_52 = 3'h4 == dispatch_io_outs_6 ? regs_4 : _GEN_51; // @[BasicChiselModules.scala 292:18]
  assign _GEN_53 = 3'h5 == dispatch_io_outs_6 ? regs_5 : _GEN_52; // @[BasicChiselModules.scala 292:18]
  assign _GEN_54 = 3'h6 == dispatch_io_outs_6 ? regs_6 : _GEN_53; // @[BasicChiselModules.scala 292:18]
  assign _GEN_55 = 3'h7 == dispatch_io_outs_6 ? regs_7 : _GEN_54; // @[BasicChiselModules.scala 292:18]
  assign _GEN_57 = 3'h1 == dispatch_io_outs_7 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_58 = 3'h2 == dispatch_io_outs_7 ? regs_2 : _GEN_57; // @[BasicChiselModules.scala 292:18]
  assign _GEN_59 = 3'h3 == dispatch_io_outs_7 ? regs_3 : _GEN_58; // @[BasicChiselModules.scala 292:18]
  assign _GEN_60 = 3'h4 == dispatch_io_outs_7 ? regs_4 : _GEN_59; // @[BasicChiselModules.scala 292:18]
  assign _GEN_61 = 3'h5 == dispatch_io_outs_7 ? regs_5 : _GEN_60; // @[BasicChiselModules.scala 292:18]
  assign _GEN_62 = 3'h6 == dispatch_io_outs_7 ? regs_6 : _GEN_61; // @[BasicChiselModules.scala 292:18]
  assign _GEN_63 = 3'h7 == dispatch_io_outs_7 ? regs_7 : _GEN_62; // @[BasicChiselModules.scala 292:18]
  assign _GEN_65 = 3'h1 == dispatch_io_outs_8 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_66 = 3'h2 == dispatch_io_outs_8 ? regs_2 : _GEN_65; // @[BasicChiselModules.scala 292:18]
  assign _GEN_67 = 3'h3 == dispatch_io_outs_8 ? regs_3 : _GEN_66; // @[BasicChiselModules.scala 292:18]
  assign _GEN_68 = 3'h4 == dispatch_io_outs_8 ? regs_4 : _GEN_67; // @[BasicChiselModules.scala 292:18]
  assign _GEN_69 = 3'h5 == dispatch_io_outs_8 ? regs_5 : _GEN_68; // @[BasicChiselModules.scala 292:18]
  assign _GEN_70 = 3'h6 == dispatch_io_outs_8 ? regs_6 : _GEN_69; // @[BasicChiselModules.scala 292:18]
  assign _GEN_71 = 3'h7 == dispatch_io_outs_8 ? regs_7 : _GEN_70; // @[BasicChiselModules.scala 292:18]
  assign _GEN_73 = 3'h1 == dispatch_io_outs_9 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_74 = 3'h2 == dispatch_io_outs_9 ? regs_2 : _GEN_73; // @[BasicChiselModules.scala 292:18]
  assign _GEN_75 = 3'h3 == dispatch_io_outs_9 ? regs_3 : _GEN_74; // @[BasicChiselModules.scala 292:18]
  assign _GEN_76 = 3'h4 == dispatch_io_outs_9 ? regs_4 : _GEN_75; // @[BasicChiselModules.scala 292:18]
  assign _GEN_77 = 3'h5 == dispatch_io_outs_9 ? regs_5 : _GEN_76; // @[BasicChiselModules.scala 292:18]
  assign _GEN_78 = 3'h6 == dispatch_io_outs_9 ? regs_6 : _GEN_77; // @[BasicChiselModules.scala 292:18]
  assign _GEN_79 = 3'h7 == dispatch_io_outs_9 ? regs_7 : _GEN_78; // @[BasicChiselModules.scala 292:18]
  assign _GEN_81 = 3'h1 == dispatch_io_outs_10 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_82 = 3'h2 == dispatch_io_outs_10 ? regs_2 : _GEN_81; // @[BasicChiselModules.scala 292:18]
  assign _GEN_83 = 3'h3 == dispatch_io_outs_10 ? regs_3 : _GEN_82; // @[BasicChiselModules.scala 292:18]
  assign _GEN_84 = 3'h4 == dispatch_io_outs_10 ? regs_4 : _GEN_83; // @[BasicChiselModules.scala 292:18]
  assign _GEN_85 = 3'h5 == dispatch_io_outs_10 ? regs_5 : _GEN_84; // @[BasicChiselModules.scala 292:18]
  assign _GEN_86 = 3'h6 == dispatch_io_outs_10 ? regs_6 : _GEN_85; // @[BasicChiselModules.scala 292:18]
  assign _GEN_87 = 3'h7 == dispatch_io_outs_10 ? regs_7 : _GEN_86; // @[BasicChiselModules.scala 292:18]
  assign _GEN_89 = 3'h1 == dispatch_io_outs_11 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_90 = 3'h2 == dispatch_io_outs_11 ? regs_2 : _GEN_89; // @[BasicChiselModules.scala 292:18]
  assign _GEN_91 = 3'h3 == dispatch_io_outs_11 ? regs_3 : _GEN_90; // @[BasicChiselModules.scala 292:18]
  assign _GEN_92 = 3'h4 == dispatch_io_outs_11 ? regs_4 : _GEN_91; // @[BasicChiselModules.scala 292:18]
  assign _GEN_93 = 3'h5 == dispatch_io_outs_11 ? regs_5 : _GEN_92; // @[BasicChiselModules.scala 292:18]
  assign _GEN_94 = 3'h6 == dispatch_io_outs_11 ? regs_6 : _GEN_93; // @[BasicChiselModules.scala 292:18]
  assign _GEN_95 = 3'h7 == dispatch_io_outs_11 ? regs_7 : _GEN_94; // @[BasicChiselModules.scala 292:18]
  assign io_outs_7 = io_en ? _GEN_95 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_6 = io_en ? _GEN_87 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_5 = io_en ? _GEN_79 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_4 = io_en ? _GEN_71 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_3 = io_en ? _GEN_63 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_2 = io_en ? _GEN_55 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_1 = io_en ? _GEN_47 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_0 = io_en ? _GEN_39 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign dispatch_io_en = io_en; // @[BasicChiselModules.scala 277:18]
  assign dispatch_io_configuration = io_configuration; // @[BasicChiselModules.scala 276:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else if (io_en) begin
      if (3'h0 == dispatch_io_outs_3) begin
        regs_0 <= io_inputs_3;
      end else if (3'h0 == dispatch_io_outs_2) begin
        regs_0 <= io_inputs_2;
      end else if (3'h0 == dispatch_io_outs_1) begin
        regs_0 <= io_inputs_1;
      end else if (3'h0 == dispatch_io_outs_0) begin
        regs_0 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_1 <= 32'h0;
    end else if (io_en) begin
      if (3'h1 == dispatch_io_outs_3) begin
        regs_1 <= io_inputs_3;
      end else if (3'h1 == dispatch_io_outs_2) begin
        regs_1 <= io_inputs_2;
      end else if (3'h1 == dispatch_io_outs_1) begin
        regs_1 <= io_inputs_1;
      end else if (3'h1 == dispatch_io_outs_0) begin
        regs_1 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'h0;
    end else if (io_en) begin
      if (3'h2 == dispatch_io_outs_3) begin
        regs_2 <= io_inputs_3;
      end else if (3'h2 == dispatch_io_outs_2) begin
        regs_2 <= io_inputs_2;
      end else if (3'h2 == dispatch_io_outs_1) begin
        regs_2 <= io_inputs_1;
      end else if (3'h2 == dispatch_io_outs_0) begin
        regs_2 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_3 <= 32'h0;
    end else if (io_en) begin
      if (3'h3 == dispatch_io_outs_3) begin
        regs_3 <= io_inputs_3;
      end else if (3'h3 == dispatch_io_outs_2) begin
        regs_3 <= io_inputs_2;
      end else if (3'h3 == dispatch_io_outs_1) begin
        regs_3 <= io_inputs_1;
      end else if (3'h3 == dispatch_io_outs_0) begin
        regs_3 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_4 <= 32'h0;
    end else if (io_en) begin
      if (3'h4 == dispatch_io_outs_3) begin
        regs_4 <= io_inputs_3;
      end else if (3'h4 == dispatch_io_outs_2) begin
        regs_4 <= io_inputs_2;
      end else if (3'h4 == dispatch_io_outs_1) begin
        regs_4 <= io_inputs_1;
      end else if (3'h4 == dispatch_io_outs_0) begin
        regs_4 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_5 <= 32'h0;
    end else if (io_en) begin
      if (3'h5 == dispatch_io_outs_3) begin
        regs_5 <= io_inputs_3;
      end else if (3'h5 == dispatch_io_outs_2) begin
        regs_5 <= io_inputs_2;
      end else if (3'h5 == dispatch_io_outs_1) begin
        regs_5 <= io_inputs_1;
      end else if (3'h5 == dispatch_io_outs_0) begin
        regs_5 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_6 <= 32'h0;
    end else if (io_en) begin
      if (3'h6 == dispatch_io_outs_3) begin
        regs_6 <= io_inputs_3;
      end else if (3'h6 == dispatch_io_outs_2) begin
        regs_6 <= io_inputs_2;
      end else if (3'h6 == dispatch_io_outs_1) begin
        regs_6 <= io_inputs_1;
      end else if (3'h6 == dispatch_io_outs_0) begin
        regs_6 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_7 <= 32'h0;
    end else if (io_en) begin
      if (3'h7 == dispatch_io_outs_3) begin
        regs_7 <= io_inputs_3;
      end else if (3'h7 == dispatch_io_outs_2) begin
        regs_7 <= io_inputs_2;
      end else if (3'h7 == dispatch_io_outs_1) begin
        regs_7 <= io_inputs_1;
      end else if (3'h7 == dispatch_io_outs_0) begin
        regs_7 <= io_inputs_0;
      end
    end
  end
endmodule
module Dispatch_2(
  input        io_en,
  input  [2:0] io_configuration,
  output       io_outs_2,
  output       io_outs_1,
  output       io_outs_0
);
  wire  _T; // @[BasicChiselModules.scala 409:37]
  wire  _T_1; // @[BasicChiselModules.scala 409:37]
  wire  _T_2; // @[BasicChiselModules.scala 409:37]
  assign _T = io_configuration[0]; // @[BasicChiselModules.scala 409:37]
  assign _T_1 = io_configuration[1]; // @[BasicChiselModules.scala 409:37]
  assign _T_2 = io_configuration[2]; // @[BasicChiselModules.scala 409:37]
  assign io_outs_2 = io_en & _T_2; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_1 = io_en & _T_1; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_0 = io_en & _T; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module RegisterFiles_1(
  input         clock,
  input         reset,
  input         io_en,
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_1,
  output [31:0] io_outs_0
);
  wire  dispatch_io_en; // @[BasicChiselModules.scala 275:24]
  wire [2:0] dispatch_io_configuration; // @[BasicChiselModules.scala 275:24]
  wire  dispatch_io_outs_2; // @[BasicChiselModules.scala 275:24]
  wire  dispatch_io_outs_1; // @[BasicChiselModules.scala 275:24]
  wire  dispatch_io_outs_0; // @[BasicChiselModules.scala 275:24]
  reg [31:0] regs_0; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[BasicChiselModules.scala 282:21]
  reg [31:0] _RAND_1;
  wire [31:0] _GEN_3; // @[BasicChiselModules.scala 292:18]
  wire [31:0] _GEN_5; // @[BasicChiselModules.scala 292:18]
  Dispatch_2 dispatch ( // @[BasicChiselModules.scala 275:24]
    .io_en(dispatch_io_en),
    .io_configuration(dispatch_io_configuration),
    .io_outs_2(dispatch_io_outs_2),
    .io_outs_1(dispatch_io_outs_1),
    .io_outs_0(dispatch_io_outs_0)
  );
  assign _GEN_3 = dispatch_io_outs_1 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign _GEN_5 = dispatch_io_outs_2 ? regs_1 : regs_0; // @[BasicChiselModules.scala 292:18]
  assign io_outs_1 = io_en ? _GEN_5 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign io_outs_0 = io_en ? _GEN_3 : 32'h0; // @[BasicChiselModules.scala 292:18 BasicChiselModules.scala 297:11]
  assign dispatch_io_en = io_en; // @[BasicChiselModules.scala 277:18]
  assign dispatch_io_configuration = io_configuration; // @[BasicChiselModules.scala 276:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'h0;
    end else if (io_en) begin
      if (1'h0 == dispatch_io_outs_0) begin
        regs_0 <= io_inputs_0;
      end
    end
    if (reset) begin
      regs_1 <= 32'h0;
    end else if (io_en) begin
      if (dispatch_io_outs_0) begin
        regs_1 <= io_inputs_0;
      end
    end
  end
endmodule
module Multiplexer(
  input         io_en,
  input  [1:0]  io_configuration,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] muxIn0; // @[Mux.scala 68:16]
  assign _T = 2'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_3 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 2'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_2 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 2'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_1 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 2'h0 == io_configuration; // @[Mux.scala 68:19]
  assign muxIn0 = _T_6 ? io_inputs_0 : _T_5; // @[Mux.scala 68:16]
  assign io_outs_0 = io_en ? muxIn0 : 32'h0; // @[BasicChiselModules.scala 317:16 BasicChiselModules.scala 320:11]
endmodule
module Multiplexer_8(
  input         io_en,
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_7,
  input  [31:0] io_inputs_6,
  input  [31:0] io_inputs_5,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  wire [31:0] _T_11; // @[Mux.scala 68:16]
  wire  _T_12; // @[Mux.scala 68:19]
  wire [31:0] _T_13; // @[Mux.scala 68:16]
  wire  _T_14; // @[Mux.scala 68:19]
  wire [31:0] muxIn0; // @[Mux.scala 68:16]
  assign _T = 3'h7 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_7 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h6 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_6 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_5 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_4 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_9 = _T_8 ? io_inputs_3 : _T_7; // @[Mux.scala 68:16]
  assign _T_10 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_11 = _T_10 ? io_inputs_2 : _T_9; // @[Mux.scala 68:16]
  assign _T_12 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_13 = _T_12 ? io_inputs_1 : _T_11; // @[Mux.scala 68:16]
  assign _T_14 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign muxIn0 = _T_14 ? io_inputs_0 : _T_13; // @[Mux.scala 68:16]
  assign io_outs_0 = io_en ? muxIn0 : 32'h0; // @[BasicChiselModules.scala 317:16 BasicChiselModules.scala 320:11]
endmodule
module Multiplexer_9(
  input         io_en,
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_6,
  input  [31:0] io_inputs_5,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  wire [31:0] _T_11; // @[Mux.scala 68:16]
  wire  _T_12; // @[Mux.scala 68:19]
  wire [31:0] muxIn0; // @[Mux.scala 68:16]
  assign _T = 3'h6 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_6 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_5 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_4 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_3 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_9 = _T_8 ? io_inputs_2 : _T_7; // @[Mux.scala 68:16]
  assign _T_10 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_11 = _T_10 ? io_inputs_1 : _T_9; // @[Mux.scala 68:16]
  assign _T_12 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign muxIn0 = _T_12 ? io_inputs_0 : _T_11; // @[Mux.scala 68:16]
  assign io_outs_0 = io_en ? muxIn0 : 32'h0; // @[BasicChiselModules.scala 317:16 BasicChiselModules.scala 320:11]
endmodule
module Multiplexer_17(
  input         io_en,
  input  [2:0]  io_configuration,
  input  [31:0] io_inputs_5,
  input  [31:0] io_inputs_4,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_0
);
  wire  _T; // @[Mux.scala 68:19]
  wire [31:0] _T_1; // @[Mux.scala 68:16]
  wire  _T_2; // @[Mux.scala 68:19]
  wire [31:0] _T_3; // @[Mux.scala 68:16]
  wire  _T_4; // @[Mux.scala 68:19]
  wire [31:0] _T_5; // @[Mux.scala 68:16]
  wire  _T_6; // @[Mux.scala 68:19]
  wire [31:0] _T_7; // @[Mux.scala 68:16]
  wire  _T_8; // @[Mux.scala 68:19]
  wire [31:0] _T_9; // @[Mux.scala 68:16]
  wire  _T_10; // @[Mux.scala 68:19]
  wire [31:0] muxIn0; // @[Mux.scala 68:16]
  assign _T = 3'h5 == io_configuration; // @[Mux.scala 68:19]
  assign _T_1 = _T ? io_inputs_5 : io_inputs_0; // @[Mux.scala 68:16]
  assign _T_2 = 3'h4 == io_configuration; // @[Mux.scala 68:19]
  assign _T_3 = _T_2 ? io_inputs_4 : _T_1; // @[Mux.scala 68:16]
  assign _T_4 = 3'h3 == io_configuration; // @[Mux.scala 68:19]
  assign _T_5 = _T_4 ? io_inputs_3 : _T_3; // @[Mux.scala 68:16]
  assign _T_6 = 3'h2 == io_configuration; // @[Mux.scala 68:19]
  assign _T_7 = _T_6 ? io_inputs_2 : _T_5; // @[Mux.scala 68:16]
  assign _T_8 = 3'h1 == io_configuration; // @[Mux.scala 68:19]
  assign _T_9 = _T_8 ? io_inputs_1 : _T_7; // @[Mux.scala 68:16]
  assign _T_10 = 3'h0 == io_configuration; // @[Mux.scala 68:19]
  assign muxIn0 = _T_10 ? io_inputs_0 : _T_9; // @[Mux.scala 68:16]
  assign io_outs_0 = io_en ? muxIn0 : 32'h0; // @[BasicChiselModules.scala 317:16 BasicChiselModules.scala 320:11]
endmodule
module ConstUnit(
  input         io_en,
  input  [31:0] io_configuration,
  output [31:0] io_outs_0
);
  assign io_outs_0 = io_en ? io_configuration : 32'h0; // @[BasicChiselModules.scala 354:16 BasicChiselModules.scala 357:11]
endmodule
module SimpleDualPortSram(
  input         clock,
  input         io_a_en,
  input         io_a_we,
  input  [7:0]  io_a_addr,
  input  [31:0] io_a_din,
  input         io_b_en,
  input  [7:0]  io_b_addr,
  output [31:0] io_b_dout
);
  reg [31:0] mem [0:255]; // @[Mem.scala 201:16]
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_2_data; // @[Mem.scala 201:16]
  wire [7:0] mem__T_2_addr; // @[Mem.scala 201:16]
  wire [31:0] mem__T_1_data; // @[Mem.scala 201:16]
  wire [7:0] mem__T_1_addr; // @[Mem.scala 201:16]
  wire  mem__T_1_mask; // @[Mem.scala 201:16]
  wire  mem__T_1_en; // @[Mem.scala 201:16]
  reg [31:0] dout; // @[Mem.scala 202:17]
  reg [31:0] _RAND_1;
  assign mem__T_2_addr = io_b_addr;
  assign mem__T_2_data = mem[mem__T_2_addr]; // @[Mem.scala 201:16]
  assign mem__T_1_data = io_a_din;
  assign mem__T_1_addr = io_a_addr;
  assign mem__T_1_mask = 1'h1;
  assign mem__T_1_en = io_a_en & io_a_we;
  assign io_b_dout = dout; // @[Mem.scala 204:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  dout = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_1_en & mem__T_1_mask) begin
      mem[mem__T_1_addr] <= mem__T_1_data; // @[Mem.scala 201:16]
    end
    if (io_b_en) begin
      dout <= mem__T_2_data;
    end
  end
endmodule
module EnqMem(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_mem_en,
  output        io_mem_we,
  output [7:0]  io_mem_addr,
  output [31:0] io_mem_din,
  input  [7:0]  io_base,
  input         io_en,
  input         io_start,
  output        io_idle
);
  reg  state; // @[EnqMem.scala 64:22]
  reg [31:0] _RAND_0;
  reg [7:0] mem_index; // @[EnqMem.scala 68:22]
  reg [31:0] _RAND_1;
  reg [31:0] data_in; // @[EnqMem.scala 69:20]
  reg [31:0] _RAND_2;
  wire  _T; // @[EnqMem.scala 75:21]
  wire  _T_1; // @[EnqMem.scala 75:38]
  wire  _T_3; // @[EnqMem.scala 79:19]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire [7:0] _T_8; // @[EnqMem.scala 95:34]
  wire  _GEN_12; // @[EnqMem.scala 91:33]
  assign _T = state == 1'h0; // @[EnqMem.scala 75:21]
  assign _T_1 = io_in_valid == 1'h0; // @[EnqMem.scala 75:38]
  assign _T_3 = io_idle & io_start; // @[EnqMem.scala 79:19]
  assign _T_5 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = mem_index + 8'h1; // @[EnqMem.scala 95:34]
  assign _GEN_12 = state | _T; // @[EnqMem.scala 91:33]
  assign io_in_ready = io_en & _GEN_12; // @[Decoupled.scala 72:20 Decoupled.scala 65:20 Decoupled.scala 65:20]
  assign io_mem_en = io_en & state; // @[Mem.scala 73:8 Mem.scala 69:8]
  assign io_mem_we = io_en & state; // @[Mem.scala 74:8 Mem.scala 70:8]
  assign io_mem_addr = mem_index; // @[EnqMem.scala 93:23]
  assign io_mem_din = data_in; // @[EnqMem.scala 94:22]
  assign io_idle = _T & _T_1; // @[EnqMem.scala 75:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_index = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  data_in = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else if (io_en) begin
      if (state) begin
        state <= _T_5;
      end else if (_T) begin
        state <= _T_5;
      end else if (_T_3) begin
        state <= 1'h0;
      end
    end
    if (io_en) begin
      if (state) begin
        mem_index <= _T_8;
      end else if (_T_3) begin
        mem_index <= io_base;
      end
    end
    if (io_en) begin
      if (state) begin
        data_in <= io_in_bits;
      end else if (_T) begin
        data_in <= io_in_bits;
      end
    end
  end
endmodule
module Handshake(
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
  assign io_enq_ready = io_deq_ready; // @[BusHelper.scala 11:10]
  assign io_deq_valid = io_enq_valid; // @[BusHelper.scala 11:10]
  assign io_deq_bits = io_enq_bits; // @[BusHelper.scala 11:10]
endmodule
module Handshake_1(
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
  assign io_enq_ready = io_deq_ready; // @[BusHelper.scala 11:10]
  assign io_deq_valid = io_enq_valid; // @[BusHelper.scala 11:10]
  assign io_deq_bits = io_enq_bits; // @[BusHelper.scala 11:10]
endmodule
module EnqAddrDeqMem(
  input         clock,
  input         reset,
  output        io_iaddr_ready,
  input         io_iaddr_valid,
  input  [7:0]  io_iaddr_bits,
  output        io_mem_en,
  output [7:0]  io_mem_addr,
  input  [31:0] io_mem_dout,
  input         io_odata_ready,
  output        io_odata_valid,
  output [31:0] io_odata_bits,
  output        io_idle
);
  reg  token; // @[DeqMem.scala 210:22]
  reg [31:0] _RAND_0;
  wire  _T; // @[DeqMem.scala 217:21]
  wire  _T_1; // @[DeqMem.scala 217:53]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_0; // @[DeqMem.scala 225:28]
  wire  _GEN_4; // @[DeqMem.scala 223:16]
  wire  _T_4; // @[DeqMem.scala 231:20]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[DeqMem.scala 233:28]
  assign _T = token == 1'h0; // @[DeqMem.scala 217:21]
  assign _T_1 = io_iaddr_valid == 1'h0; // @[DeqMem.scala 217:53]
  assign _T_3 = io_odata_ready & io_odata_valid; // @[Decoupled.scala 40:37]
  assign _GEN_0 = _T_3 ? 1'h0 : token; // @[DeqMem.scala 225:28]
  assign _GEN_4 = token ? _GEN_0 : token; // @[DeqMem.scala 223:16]
  assign _T_4 = _GEN_4 == 1'h0; // @[DeqMem.scala 231:20]
  assign _T_5 = io_iaddr_ready & io_iaddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_5 | _GEN_4; // @[DeqMem.scala 233:28]
  assign io_iaddr_ready = _GEN_4 == 1'h0; // @[Decoupled.scala 72:20 Decoupled.scala 65:20]
  assign io_mem_en = _T_4 & _T_5; // @[Mem.scala 43:8 Mem.scala 40:8]
  assign io_mem_addr = io_iaddr_bits; // @[DeqMem.scala 236:19]
  assign io_odata_valid = token; // @[Decoupled.scala 56:20 Decoupled.scala 47:20]
  assign io_odata_bits = io_mem_dout; // @[Decoupled.scala 48:19]
  assign io_idle = _T & _T_1; // @[DeqMem.scala 217:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  token = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      token <= 1'h0;
    end else if (_T_4) begin
      token <= _GEN_6;
    end else if (token) begin
      if (_T_3) begin
        token <= 1'h0;
      end
    end
  end
endmodule
module DeqMem(
  input         clock,
  input         reset,
  output        io_mem_en,
  output [7:0]  io_mem_addr,
  input  [31:0] io_mem_dout,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits,
  input  [7:0]  io_base,
  input  [7:0]  io_len,
  input         io_en,
  input         io_start,
  output        io_idle
);
  wire  iaddr_hs_io_enq_ready; // @[DeqMem.scala 100:24]
  wire  iaddr_hs_io_enq_valid; // @[DeqMem.scala 100:24]
  wire [7:0] iaddr_hs_io_enq_bits; // @[DeqMem.scala 100:24]
  wire  iaddr_hs_io_deq_ready; // @[DeqMem.scala 100:24]
  wire  iaddr_hs_io_deq_valid; // @[DeqMem.scala 100:24]
  wire [7:0] iaddr_hs_io_deq_bits; // @[DeqMem.scala 100:24]
  wire  odata_hs_io_enq_ready; // @[DeqMem.scala 103:24]
  wire  odata_hs_io_enq_valid; // @[DeqMem.scala 103:24]
  wire [31:0] odata_hs_io_enq_bits; // @[DeqMem.scala 103:24]
  wire  odata_hs_io_deq_ready; // @[DeqMem.scala 103:24]
  wire  odata_hs_io_deq_valid; // @[DeqMem.scala 103:24]
  wire [31:0] odata_hs_io_deq_bits; // @[DeqMem.scala 103:24]
  wire  EnqAddrDeqMem_clock; // @[DeqMem.scala 54:22]
  wire  EnqAddrDeqMem_reset; // @[DeqMem.scala 54:22]
  wire  EnqAddrDeqMem_io_iaddr_ready; // @[DeqMem.scala 54:22]
  wire  EnqAddrDeqMem_io_iaddr_valid; // @[DeqMem.scala 54:22]
  wire [7:0] EnqAddrDeqMem_io_iaddr_bits; // @[DeqMem.scala 54:22]
  wire  EnqAddrDeqMem_io_mem_en; // @[DeqMem.scala 54:22]
  wire [7:0] EnqAddrDeqMem_io_mem_addr; // @[DeqMem.scala 54:22]
  wire [31:0] EnqAddrDeqMem_io_mem_dout; // @[DeqMem.scala 54:22]
  wire  EnqAddrDeqMem_io_odata_ready; // @[DeqMem.scala 54:22]
  wire  EnqAddrDeqMem_io_odata_valid; // @[DeqMem.scala 54:22]
  wire [31:0] EnqAddrDeqMem_io_odata_bits; // @[DeqMem.scala 54:22]
  wire  EnqAddrDeqMem_io_idle; // @[DeqMem.scala 54:22]
  reg [1:0] state; // @[DeqMem.scala 91:22]
  reg [31:0] _RAND_0;
  reg [7:0] mem_index; // @[DeqMem.scala 95:22]
  reg [31:0] _RAND_1;
  reg [31:0] mem_data; // @[DeqMem.scala 96:21]
  reg [31:0] _RAND_2;
  reg [7:0] remain; // @[DeqMem.scala 98:19]
  reg [31:0] _RAND_3;
  wire  _T_1; // @[DeqMem.scala 121:19]
  wire [7:0] _GEN_1; // @[DeqMem.scala 121:32]
  wire [7:0] _GEN_3; // @[DeqMem.scala 121:32]
  wire  _T_2; // @[DeqMem.scala 128:17]
  wire  _T_3; // @[DeqMem.scala 183:18]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire [7:0] _T_6; // @[DeqMem.scala 186:32]
  wire [7:0] _T_8; // @[DeqMem.scala 187:26]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[DeqMem.scala 194:29]
  wire  _GEN_12; // @[DeqMem.scala 128:30]
  wire  _T_11; // @[DeqMem.scala 134:21]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[DeqMem.scala 183:25]
  wire  _GEN_27; // @[DeqMem.scala 136:32]
  wire  _GEN_31; // @[DeqMem.scala 136:32]
  wire  _GEN_36; // @[DeqMem.scala 134:33]
  wire  _GEN_40; // @[DeqMem.scala 134:33]
  Handshake iaddr_hs ( // @[DeqMem.scala 100:24]
    .io_enq_ready(iaddr_hs_io_enq_ready),
    .io_enq_valid(iaddr_hs_io_enq_valid),
    .io_enq_bits(iaddr_hs_io_enq_bits),
    .io_deq_ready(iaddr_hs_io_deq_ready),
    .io_deq_valid(iaddr_hs_io_deq_valid),
    .io_deq_bits(iaddr_hs_io_deq_bits)
  );
  Handshake_1 odata_hs ( // @[DeqMem.scala 103:24]
    .io_enq_ready(odata_hs_io_enq_ready),
    .io_enq_valid(odata_hs_io_enq_valid),
    .io_enq_bits(odata_hs_io_enq_bits),
    .io_deq_ready(odata_hs_io_deq_ready),
    .io_deq_valid(odata_hs_io_deq_valid),
    .io_deq_bits(odata_hs_io_deq_bits)
  );
  EnqAddrDeqMem EnqAddrDeqMem ( // @[DeqMem.scala 54:22]
    .clock(EnqAddrDeqMem_clock),
    .reset(EnqAddrDeqMem_reset),
    .io_iaddr_ready(EnqAddrDeqMem_io_iaddr_ready),
    .io_iaddr_valid(EnqAddrDeqMem_io_iaddr_valid),
    .io_iaddr_bits(EnqAddrDeqMem_io_iaddr_bits),
    .io_mem_en(EnqAddrDeqMem_io_mem_en),
    .io_mem_addr(EnqAddrDeqMem_io_mem_addr),
    .io_mem_dout(EnqAddrDeqMem_io_mem_dout),
    .io_odata_ready(EnqAddrDeqMem_io_odata_ready),
    .io_odata_valid(EnqAddrDeqMem_io_odata_valid),
    .io_odata_bits(EnqAddrDeqMem_io_odata_bits),
    .io_idle(EnqAddrDeqMem_io_idle)
  );
  assign _T_1 = io_idle & io_start; // @[DeqMem.scala 121:19]
  assign _GEN_1 = _T_1 ? io_base : mem_index; // @[DeqMem.scala 121:32]
  assign _GEN_3 = _T_1 ? io_len : remain; // @[DeqMem.scala 121:32]
  assign _T_2 = state == 2'h1; // @[DeqMem.scala 128:17]
  assign _T_3 = remain > 8'h0; // @[DeqMem.scala 183:18]
  assign _T_4 = iaddr_hs_io_enq_ready & iaddr_hs_io_enq_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = mem_index + 8'h1; // @[DeqMem.scala 186:32]
  assign _T_8 = remain - 8'h1; // @[DeqMem.scala 187:26]
  assign _T_9 = odata_hs_io_deq_ready & odata_hs_io_deq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = EnqAddrDeqMem_io_idle == 1'h0; // @[DeqMem.scala 194:29]
  assign _GEN_12 = _T_2 & _T_3; // @[DeqMem.scala 128:30]
  assign _T_11 = state == 2'h2; // @[DeqMem.scala 134:21]
  assign _T_12 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_3 | _GEN_12; // @[DeqMem.scala 183:25]
  assign _GEN_27 = _T_12 ? _GEN_21 : _GEN_12; // @[DeqMem.scala 136:32]
  assign _GEN_31 = _T_12 | _T_2; // @[DeqMem.scala 136:32]
  assign _GEN_36 = _T_11 ? _GEN_27 : _GEN_12; // @[DeqMem.scala 134:33]
  assign _GEN_40 = _T_11 ? _GEN_31 : _T_2; // @[DeqMem.scala 134:33]
  assign io_mem_en = EnqAddrDeqMem_io_mem_en; // @[Mem.scala 43:8 DeqMem.scala 68:22]
  assign io_mem_addr = EnqAddrDeqMem_io_mem_addr; // @[DeqMem.scala 69:24]
  assign io_out_valid = io_en & _T_11; // @[Decoupled.scala 56:20 Decoupled.scala 47:20]
  assign io_out_bits = mem_data; // @[Decoupled.scala 48:19]
  assign io_idle = state == 2'h0; // @[DeqMem.scala 115:11]
  assign iaddr_hs_io_enq_valid = io_en & _GEN_36; // @[Decoupled.scala 56:20 Decoupled.scala 47:20 Decoupled.scala 47:20]
  assign iaddr_hs_io_enq_bits = mem_index; // @[Decoupled.scala 48:19 Decoupled.scala 48:19]
  assign iaddr_hs_io_deq_ready = EnqAddrDeqMem_io_iaddr_ready; // @[Decoupled.scala 72:20 DeqMem.scala 67:21]
  assign odata_hs_io_enq_valid = EnqAddrDeqMem_io_odata_valid; // @[Decoupled.scala 56:20 DeqMem.scala 71:21]
  assign odata_hs_io_enq_bits = EnqAddrDeqMem_io_odata_bits; // @[DeqMem.scala 71:21]
  assign odata_hs_io_deq_ready = io_en & _GEN_40; // @[Decoupled.scala 72:20 Decoupled.scala 65:20 Decoupled.scala 65:20]
  assign EnqAddrDeqMem_clock = clock;
  assign EnqAddrDeqMem_reset = reset;
  assign EnqAddrDeqMem_io_iaddr_valid = iaddr_hs_io_deq_valid; // @[Decoupled.scala 56:20 DeqMem.scala 67:21]
  assign EnqAddrDeqMem_io_iaddr_bits = iaddr_hs_io_deq_bits; // @[DeqMem.scala 67:21]
  assign EnqAddrDeqMem_io_mem_dout = io_mem_dout; // @[DeqMem.scala 70:24]
  assign EnqAddrDeqMem_io_odata_ready = odata_hs_io_enq_ready; // @[Decoupled.scala 72:20 DeqMem.scala 71:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_index = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  remain = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          if (_T_9) begin
            state <= 2'h2;
          end else if (_T_10) begin
            state <= 2'h1;
          end else begin
            state <= 2'h0;
          end
        end else if (_T_2) begin
          if (_T_9) begin
            state <= 2'h2;
          end else if (_T_10) begin
            state <= 2'h1;
          end else begin
            state <= 2'h0;
          end
        end else if (_T_1) begin
          state <= 2'h1;
        end
      end else if (_T_2) begin
        if (_T_9) begin
          state <= 2'h2;
        end else if (_T_10) begin
          state <= 2'h1;
        end else begin
          state <= 2'h0;
        end
      end else if (_T_1) begin
        state <= 2'h1;
      end
    end
    if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          if (_T_3) begin
            if (_T_4) begin
              mem_index <= _T_6;
            end else if (_T_2) begin
              if (_T_3) begin
                if (_T_4) begin
                  mem_index <= _T_6;
                end else if (_T_1) begin
                  mem_index <= io_base;
                end
              end else if (_T_1) begin
                mem_index <= io_base;
              end
            end else if (_T_1) begin
              mem_index <= io_base;
            end
          end else if (_T_2) begin
            if (_T_3) begin
              if (_T_4) begin
                mem_index <= _T_6;
              end else if (_T_1) begin
                mem_index <= io_base;
              end
            end else begin
              mem_index <= _GEN_1;
            end
          end else begin
            mem_index <= _GEN_1;
          end
        end else if (_T_2) begin
          if (_T_3) begin
            if (_T_4) begin
              mem_index <= _T_6;
            end else begin
              mem_index <= _GEN_1;
            end
          end else begin
            mem_index <= _GEN_1;
          end
        end else begin
          mem_index <= _GEN_1;
        end
      end else if (_T_2) begin
        if (_T_3) begin
          if (_T_4) begin
            mem_index <= _T_6;
          end else begin
            mem_index <= _GEN_1;
          end
        end else begin
          mem_index <= _GEN_1;
        end
      end else begin
        mem_index <= _GEN_1;
      end
    end
    if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          mem_data <= odata_hs_io_deq_bits;
        end else if (_T_2) begin
          mem_data <= odata_hs_io_deq_bits;
        end
      end else if (_T_2) begin
        mem_data <= odata_hs_io_deq_bits;
      end
    end
    if (io_en) begin
      if (_T_11) begin
        if (_T_12) begin
          if (_T_3) begin
            if (_T_4) begin
              remain <= _T_8;
            end else if (_T_2) begin
              if (_T_3) begin
                if (_T_4) begin
                  remain <= _T_8;
                end else if (_T_1) begin
                  remain <= io_len;
                end
              end else if (_T_1) begin
                remain <= io_len;
              end
            end else if (_T_1) begin
              remain <= io_len;
            end
          end else if (_T_2) begin
            if (_T_3) begin
              if (_T_4) begin
                remain <= _T_8;
              end else if (_T_1) begin
                remain <= io_len;
              end
            end else begin
              remain <= _GEN_3;
            end
          end else begin
            remain <= _GEN_3;
          end
        end else if (_T_2) begin
          if (_T_3) begin
            if (_T_4) begin
              remain <= _T_8;
            end else begin
              remain <= _GEN_3;
            end
          end else begin
            remain <= _GEN_3;
          end
        end else begin
          remain <= _GEN_3;
        end
      end else if (_T_2) begin
        if (_T_3) begin
          if (_T_4) begin
            remain <= _T_8;
          end else begin
            remain <= _GEN_3;
          end
        end else begin
          remain <= _GEN_3;
        end
      end else begin
        remain <= _GEN_3;
      end
    end
  end
endmodule
module LSMemWrapper(
  input         clock,
  input         reset,
  input         io_workEn,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  input         io_readMem_en,
  input  [7:0]  io_readMem_addr,
  output [31:0] io_readMem_dout,
  input         io_writeMem_en,
  input         io_writeMem_we,
  input  [7:0]  io_writeMem_addr,
  input  [31:0] io_writeMem_din,
  input  [7:0]  io_base,
  input  [7:0]  io_len,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits,
  input         io_start,
  input         io_enqEn,
  input         io_deqEn,
  output        io_idle
);
  wire  mem_clock; // @[BasicChiselModules.scala 459:19]
  wire  mem_io_a_en; // @[BasicChiselModules.scala 459:19]
  wire  mem_io_a_we; // @[BasicChiselModules.scala 459:19]
  wire [7:0] mem_io_a_addr; // @[BasicChiselModules.scala 459:19]
  wire [31:0] mem_io_a_din; // @[BasicChiselModules.scala 459:19]
  wire  mem_io_b_en; // @[BasicChiselModules.scala 459:19]
  wire [7:0] mem_io_b_addr; // @[BasicChiselModules.scala 459:19]
  wire [31:0] mem_io_b_dout; // @[BasicChiselModules.scala 459:19]
  wire  enq_mem_clock; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_reset; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_io_in_ready; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_io_in_valid; // @[BasicChiselModules.scala 460:23]
  wire [31:0] enq_mem_io_in_bits; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_io_mem_en; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_io_mem_we; // @[BasicChiselModules.scala 460:23]
  wire [7:0] enq_mem_io_mem_addr; // @[BasicChiselModules.scala 460:23]
  wire [31:0] enq_mem_io_mem_din; // @[BasicChiselModules.scala 460:23]
  wire [7:0] enq_mem_io_base; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_io_en; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_io_start; // @[BasicChiselModules.scala 460:23]
  wire  enq_mem_io_idle; // @[BasicChiselModules.scala 460:23]
  wire  deq_mem_clock; // @[BasicChiselModules.scala 461:23]
  wire  deq_mem_reset; // @[BasicChiselModules.scala 461:23]
  wire  deq_mem_io_mem_en; // @[BasicChiselModules.scala 461:23]
  wire [7:0] deq_mem_io_mem_addr; // @[BasicChiselModules.scala 461:23]
  wire [31:0] deq_mem_io_mem_dout; // @[BasicChiselModules.scala 461:23]
  wire  deq_mem_io_out_ready; // @[BasicChiselModules.scala 461:23]
  wire  deq_mem_io_out_valid; // @[BasicChiselModules.scala 461:23]
  wire [31:0] deq_mem_io_out_bits; // @[BasicChiselModules.scala 461:23]
  wire [7:0] deq_mem_io_base; // @[BasicChiselModules.scala 461:23]
  wire [7:0] deq_mem_io_len; // @[BasicChiselModules.scala 461:23]
  wire  deq_mem_io_en; // @[BasicChiselModules.scala 461:23]
  wire  deq_mem_io_start; // @[BasicChiselModules.scala 461:23]
  wire  deq_mem_io_idle; // @[BasicChiselModules.scala 461:23]
  reg [1:0] state; // @[BasicChiselModules.scala 457:22]
  reg [31:0] _RAND_0;
  wire  _T; // @[BasicChiselModules.scala 463:14]
  wire  _GEN_1; // @[BasicChiselModules.scala 468:32]
  wire  _GEN_2; // @[BasicChiselModules.scala 468:32]
  wire [7:0] _GEN_3; // @[BasicChiselModules.scala 468:32]
  wire [31:0] _GEN_4; // @[BasicChiselModules.scala 468:32]
  wire  _GEN_6; // @[BasicChiselModules.scala 464:31]
  wire  _GEN_7; // @[BasicChiselModules.scala 464:31]
  wire [7:0] _GEN_8; // @[BasicChiselModules.scala 464:31]
  wire [31:0] _GEN_9; // @[BasicChiselModules.scala 464:31]
  wire  _T_3; // @[BasicChiselModules.scala 478:20]
  wire  _T_4; // @[BasicChiselModules.scala 479:19]
  wire  _GEN_11; // @[BasicChiselModules.scala 479:31]
  wire  _GEN_12; // @[BasicChiselModules.scala 479:31]
  wire [7:0] _GEN_13; // @[BasicChiselModules.scala 479:31]
  wire [31:0] _GEN_14; // @[BasicChiselModules.scala 479:31]
  wire  _T_5; // @[BasicChiselModules.scala 488:20]
  wire  _GEN_16; // @[BasicChiselModules.scala 489:30]
  wire [7:0] _GEN_17; // @[BasicChiselModules.scala 489:30]
  wire [31:0] _GEN_18; // @[BasicChiselModules.scala 489:30]
  wire  _T_7; // @[BasicChiselModules.scala 500:19]
  wire  _GEN_21; // @[BasicChiselModules.scala 500:31]
  wire [7:0] _GEN_22; // @[BasicChiselModules.scala 500:31]
  wire  _GEN_26; // @[BasicChiselModules.scala 488:31]
  wire [7:0] _GEN_27; // @[BasicChiselModules.scala 488:31]
  wire [31:0] _GEN_28; // @[BasicChiselModules.scala 488:31]
  wire  _GEN_34; // @[BasicChiselModules.scala 488:31]
  wire  _GEN_36; // @[BasicChiselModules.scala 478:38]
  wire  _GEN_37; // @[BasicChiselModules.scala 478:38]
  wire [7:0] _GEN_38; // @[BasicChiselModules.scala 478:38]
  wire [31:0] _GEN_39; // @[BasicChiselModules.scala 478:38]
  wire  _GEN_40; // @[BasicChiselModules.scala 478:38]
  wire [7:0] _GEN_41; // @[BasicChiselModules.scala 478:38]
  wire [31:0] _GEN_42; // @[BasicChiselModules.scala 478:38]
  wire  _GEN_44; // @[BasicChiselModules.scala 478:38]
  SimpleDualPortSram mem ( // @[BasicChiselModules.scala 459:19]
    .clock(mem_clock),
    .io_a_en(mem_io_a_en),
    .io_a_we(mem_io_a_we),
    .io_a_addr(mem_io_a_addr),
    .io_a_din(mem_io_a_din),
    .io_b_en(mem_io_b_en),
    .io_b_addr(mem_io_b_addr),
    .io_b_dout(mem_io_b_dout)
  );
  EnqMem enq_mem ( // @[BasicChiselModules.scala 460:23]
    .clock(enq_mem_clock),
    .reset(enq_mem_reset),
    .io_in_ready(enq_mem_io_in_ready),
    .io_in_valid(enq_mem_io_in_valid),
    .io_in_bits(enq_mem_io_in_bits),
    .io_mem_en(enq_mem_io_mem_en),
    .io_mem_we(enq_mem_io_mem_we),
    .io_mem_addr(enq_mem_io_mem_addr),
    .io_mem_din(enq_mem_io_mem_din),
    .io_base(enq_mem_io_base),
    .io_en(enq_mem_io_en),
    .io_start(enq_mem_io_start),
    .io_idle(enq_mem_io_idle)
  );
  DeqMem deq_mem ( // @[BasicChiselModules.scala 461:23]
    .clock(deq_mem_clock),
    .reset(deq_mem_reset),
    .io_mem_en(deq_mem_io_mem_en),
    .io_mem_addr(deq_mem_io_mem_addr),
    .io_mem_dout(deq_mem_io_mem_dout),
    .io_out_ready(deq_mem_io_out_ready),
    .io_out_valid(deq_mem_io_out_valid),
    .io_out_bits(deq_mem_io_out_bits),
    .io_base(deq_mem_io_base),
    .io_len(deq_mem_io_len),
    .io_en(deq_mem_io_en),
    .io_start(deq_mem_io_start),
    .io_idle(deq_mem_io_idle)
  );
  assign _T = state == 2'h0; // @[BasicChiselModules.scala 463:14]
  assign _GEN_1 = io_enqEn ? enq_mem_io_mem_en : io_writeMem_en; // @[BasicChiselModules.scala 468:32]
  assign _GEN_2 = io_enqEn ? enq_mem_io_mem_we : io_writeMem_we; // @[BasicChiselModules.scala 468:32]
  assign _GEN_3 = io_enqEn ? enq_mem_io_mem_addr : io_writeMem_addr; // @[BasicChiselModules.scala 468:32]
  assign _GEN_4 = io_enqEn ? enq_mem_io_mem_din : io_writeMem_din; // @[BasicChiselModules.scala 468:32]
  assign _GEN_6 = io_workEn ? io_writeMem_en : _GEN_1; // @[BasicChiselModules.scala 464:31]
  assign _GEN_7 = io_workEn ? io_writeMem_we : _GEN_2; // @[BasicChiselModules.scala 464:31]
  assign _GEN_8 = io_workEn ? io_writeMem_addr : _GEN_3; // @[BasicChiselModules.scala 464:31]
  assign _GEN_9 = io_workEn ? io_writeMem_din : _GEN_4; // @[BasicChiselModules.scala 464:31]
  assign _T_3 = state == 2'h1; // @[BasicChiselModules.scala 478:20]
  assign _T_4 = io_enqEn == 1'h0; // @[BasicChiselModules.scala 479:19]
  assign _GEN_11 = _T_4 ? io_writeMem_en : enq_mem_io_mem_en; // @[BasicChiselModules.scala 479:31]
  assign _GEN_12 = _T_4 ? io_writeMem_we : enq_mem_io_mem_we; // @[BasicChiselModules.scala 479:31]
  assign _GEN_13 = _T_4 ? io_writeMem_addr : enq_mem_io_mem_addr; // @[BasicChiselModules.scala 479:31]
  assign _GEN_14 = _T_4 ? io_writeMem_din : enq_mem_io_mem_din; // @[BasicChiselModules.scala 479:31]
  assign _T_5 = state == 2'h2; // @[BasicChiselModules.scala 488:20]
  assign _GEN_16 = io_deqEn ? deq_mem_io_mem_en : io_readMem_en; // @[BasicChiselModules.scala 489:30]
  assign _GEN_17 = io_deqEn ? deq_mem_io_mem_addr : io_readMem_addr; // @[BasicChiselModules.scala 489:30]
  assign _GEN_18 = mem_io_b_dout; // @[BasicChiselModules.scala 489:30]
  assign _T_7 = io_deqEn == 1'h0; // @[BasicChiselModules.scala 500:19]
  assign _GEN_21 = _T_7 ? io_readMem_en : deq_mem_io_mem_en; // @[BasicChiselModules.scala 500:31]
  assign _GEN_22 = _T_7 ? io_readMem_addr : deq_mem_io_mem_addr; // @[BasicChiselModules.scala 500:31]
  assign _GEN_26 = _T_5 ? _GEN_16 : _GEN_21; // @[BasicChiselModules.scala 488:31]
  assign _GEN_27 = _T_5 ? _GEN_17 : _GEN_22; // @[BasicChiselModules.scala 488:31]
  assign _GEN_28 = _T_5 ? _GEN_18 : _GEN_18; // @[BasicChiselModules.scala 488:31]
  assign _GEN_34 = deq_mem_io_idle; // @[BasicChiselModules.scala 488:31]
  assign _GEN_36 = _T_3 ? _GEN_11 : io_writeMem_en; // @[BasicChiselModules.scala 478:38]
  assign _GEN_37 = _T_3 ? _GEN_12 : io_writeMem_we; // @[BasicChiselModules.scala 478:38]
  assign _GEN_38 = _T_3 ? _GEN_13 : io_writeMem_addr; // @[BasicChiselModules.scala 478:38]
  assign _GEN_39 = _T_3 ? _GEN_14 : io_writeMem_din; // @[BasicChiselModules.scala 478:38]
  assign _GEN_40 = _T_3 ? io_readMem_en : _GEN_26; // @[BasicChiselModules.scala 478:38]
  assign _GEN_41 = _T_3 ? io_readMem_addr : _GEN_27; // @[BasicChiselModules.scala 478:38]
  assign _GEN_42 = _T_3 ? mem_io_b_dout : _GEN_28; // @[BasicChiselModules.scala 478:38]
  assign _GEN_44 = _T_3 ? enq_mem_io_idle : _GEN_34; // @[BasicChiselModules.scala 478:38]
  assign io_in_ready = enq_mem_io_in_ready; // @[BasicChiselModules.scala 536:17]
  assign io_readMem_dout = _T ? mem_io_b_dout : _GEN_42; // @[Mem.scala 55:15 Mem.scala 55:15 Mem.scala 55:15 Mem.scala 55:15]
  assign io_out_valid = deq_mem_io_out_valid; // @[BasicChiselModules.scala 540:18]
  assign io_out_bits = deq_mem_io_out_bits; // @[BasicChiselModules.scala 540:18]
  assign io_idle = _T ? enq_mem_io_idle : _GEN_44; // @[BasicChiselModules.scala 477:21 BasicChiselModules.scala 487:21 BasicChiselModules.scala 498:21 BasicChiselModules.scala 509:21]
  assign mem_clock = clock; // @[BasicChiselModules.scala 520:13]
  assign mem_io_a_en = _T ? _GEN_6 : _GEN_36; // @[Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13 Mem.scala 90:13]
  assign mem_io_a_we = _T ? _GEN_7 : _GEN_37; // @[Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13 Mem.scala 91:13]
  assign mem_io_a_addr = _T ? _GEN_8 : _GEN_38; // @[Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15 Mem.scala 92:15]
  assign mem_io_a_din = _T ? _GEN_9 : _GEN_39; // @[Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14 Mem.scala 93:14]
  assign mem_io_b_en = _T ? io_readMem_en : _GEN_40; // @[Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13 Mem.scala 53:13]
  assign mem_io_b_addr = _T ? io_readMem_addr : _GEN_41; // @[Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15 Mem.scala 54:15]
  assign enq_mem_clock = clock; // @[BasicChiselModules.scala 521:17]
  assign enq_mem_reset = reset;
  assign enq_mem_io_in_valid = io_in_valid; // @[BasicChiselModules.scala 536:17]
  assign enq_mem_io_in_bits = io_in_bits; // @[BasicChiselModules.scala 536:17]
  assign enq_mem_io_base = io_base; // @[BasicChiselModules.scala 525:19]
  assign enq_mem_io_en = io_enqEn; // @[BasicChiselModules.scala 535:17]
  assign enq_mem_io_start = io_start; // @[BasicChiselModules.scala 526:20]
  assign deq_mem_clock = clock;
  assign deq_mem_reset = reset;
  assign deq_mem_io_mem_dout = _T_5 ? _GEN_18 : _GEN_18; // @[Mem.scala 55:15 Mem.scala 55:15]
  assign deq_mem_io_out_ready = io_out_ready; // @[BasicChiselModules.scala 540:18]
  assign deq_mem_io_base = io_base; // @[BasicChiselModules.scala 523:19]
  assign deq_mem_io_len = io_len; // @[BasicChiselModules.scala 539:18]
  assign deq_mem_io_en = io_deqEn; // @[BasicChiselModules.scala 538:17]
  assign deq_mem_io_start = io_start; // @[BasicChiselModules.scala 524:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T) begin
      if (io_workEn) begin
        state <= 2'h2;
      end else if (io_enqEn) begin
        state <= 2'h1;
      end
    end else if (_T_3) begin
      if (_T_4) begin
        state <= 2'h2;
      end
    end else if (_T_5) begin
      if (io_deqEn) begin
        state <= 2'h3;
      end
    end else if (_T_7) begin
      state <= 2'h0;
    end
  end
endmodule
module LoadStoreUnit(
  input         clock,
  input         reset,
  input         io_configuration,
  input         io_en,
  input  [4:0]  io_skewing,
  output        io_streamIn_ready,
  input         io_streamIn_valid,
  input  [31:0] io_streamIn_bits,
  input  [7:0]  io_len,
  input         io_streamOut_ready,
  output        io_streamOut_valid,
  output [31:0] io_streamOut_bits,
  input  [7:0]  io_base,
  input         io_start,
  input         io_enqEn,
  input         io_deqEn,
  output        io_idle,
  input  [31:0] io_inputs_1,
  input  [7:0]  io_inputs_0,
  output [31:0] io_outs_0
);
  wire  memWrapper_clock; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_reset; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_workEn; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_in_ready; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_in_valid; // @[BasicChiselModules.scala 567:26]
  wire [31:0] memWrapper_io_in_bits; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_readMem_en; // @[BasicChiselModules.scala 567:26]
  wire [7:0] memWrapper_io_readMem_addr; // @[BasicChiselModules.scala 567:26]
  wire [31:0] memWrapper_io_readMem_dout; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_writeMem_en; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_writeMem_we; // @[BasicChiselModules.scala 567:26]
  wire [7:0] memWrapper_io_writeMem_addr; // @[BasicChiselModules.scala 567:26]
  wire [31:0] memWrapper_io_writeMem_din; // @[BasicChiselModules.scala 567:26]
  wire [7:0] memWrapper_io_base; // @[BasicChiselModules.scala 567:26]
  wire [7:0] memWrapper_io_len; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_out_ready; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_out_valid; // @[BasicChiselModules.scala 567:26]
  wire [31:0] memWrapper_io_out_bits; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_start; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_enqEn; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_deqEn; // @[BasicChiselModules.scala 567:26]
  wire  memWrapper_io_idle; // @[BasicChiselModules.scala 567:26]
  wire  syncScheduleController_clock; // @[BasicChiselModules.scala 578:38]
  wire  syncScheduleController_reset; // @[BasicChiselModules.scala 578:38]
  wire [4:0] syncScheduleController_io_skewing; // @[BasicChiselModules.scala 578:38]
  wire [31:0] syncScheduleController_io_input0; // @[BasicChiselModules.scala 578:38]
  wire [31:0] syncScheduleController_io_input1; // @[BasicChiselModules.scala 578:38]
  wire [31:0] syncScheduleController_io_skewedInput0; // @[BasicChiselModules.scala 578:38]
  wire [31:0] syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 578:38]
  wire  _T; // @[BasicChiselModules.scala 597:27]
  wire  _GEN_1; // @[BasicChiselModules.scala 597:35]
  wire [31:0] _GEN_2; // @[BasicChiselModules.scala 593:14]
  LSMemWrapper memWrapper ( // @[BasicChiselModules.scala 567:26]
    .clock(memWrapper_clock),
    .reset(memWrapper_reset),
    .io_workEn(memWrapper_io_workEn),
    .io_in_ready(memWrapper_io_in_ready),
    .io_in_valid(memWrapper_io_in_valid),
    .io_in_bits(memWrapper_io_in_bits),
    .io_readMem_en(memWrapper_io_readMem_en),
    .io_readMem_addr(memWrapper_io_readMem_addr),
    .io_readMem_dout(memWrapper_io_readMem_dout),
    .io_writeMem_en(memWrapper_io_writeMem_en),
    .io_writeMem_we(memWrapper_io_writeMem_we),
    .io_writeMem_addr(memWrapper_io_writeMem_addr),
    .io_writeMem_din(memWrapper_io_writeMem_din),
    .io_base(memWrapper_io_base),
    .io_len(memWrapper_io_len),
    .io_out_ready(memWrapper_io_out_ready),
    .io_out_valid(memWrapper_io_out_valid),
    .io_out_bits(memWrapper_io_out_bits),
    .io_start(memWrapper_io_start),
    .io_enqEn(memWrapper_io_enqEn),
    .io_deqEn(memWrapper_io_deqEn),
    .io_idle(memWrapper_io_idle)
  );
  SyncScheduleController syncScheduleController ( // @[BasicChiselModules.scala 578:38]
    .clock(syncScheduleController_clock),
    .reset(syncScheduleController_reset),
    .io_skewing(syncScheduleController_io_skewing),
    .io_input0(syncScheduleController_io_input0),
    .io_input1(syncScheduleController_io_input1),
    .io_skewedInput0(syncScheduleController_io_skewedInput0),
    .io_skewedInput1(syncScheduleController_io_skewedInput1)
  );
  assign _T = io_configuration == 1'h0; // @[BasicChiselModules.scala 597:27]
  assign _GEN_1 = _T ? 1'h0 : 1'h1; // @[BasicChiselModules.scala 597:35]
  assign _GEN_2 = syncScheduleController_io_skewedInput0; // @[BasicChiselModules.scala 593:14]
  assign io_streamIn_ready = memWrapper_io_in_ready; // @[BasicChiselModules.scala 574:20]
  assign io_streamOut_valid = memWrapper_io_out_valid; // @[BasicChiselModules.scala 575:21]
  assign io_streamOut_bits = memWrapper_io_out_bits; // @[BasicChiselModules.scala 575:21]
  assign io_idle = memWrapper_io_idle; // @[BasicChiselModules.scala 570:22]
  assign io_outs_0 = io_en ? memWrapper_io_readMem_dout : 32'h0; // @[BasicChiselModules.scala 606:16 BasicChiselModules.scala 615:13]
  assign memWrapper_clock = clock;
  assign memWrapper_reset = reset;
  assign memWrapper_io_workEn = io_en; // @[BasicChiselModules.scala 576:24]
  assign memWrapper_io_in_valid = io_streamIn_valid; // @[BasicChiselModules.scala 574:20]
  assign memWrapper_io_in_bits = io_streamIn_bits; // @[BasicChiselModules.scala 574:20]
  assign memWrapper_io_readMem_en = io_en & _T; // @[BasicChiselModules.scala 598:18 BasicChiselModules.scala 602:18 BasicChiselModules.scala 608:16]
  assign memWrapper_io_readMem_addr = _GEN_2[7:0]; // @[BasicChiselModules.scala 594:18]
  assign memWrapper_io_writeMem_en = io_en & _GEN_1; // @[BasicChiselModules.scala 599:19 BasicChiselModules.scala 603:19 BasicChiselModules.scala 609:17]
  assign memWrapper_io_writeMem_we = io_en & _GEN_1; // @[BasicChiselModules.scala 600:19 BasicChiselModules.scala 604:19 BasicChiselModules.scala 610:17]
  assign memWrapper_io_writeMem_addr = _GEN_2[7:0]; // @[BasicChiselModules.scala 595:19]
  assign memWrapper_io_writeMem_din = syncScheduleController_io_skewedInput1; // @[BasicChiselModules.scala 596:18]
  assign memWrapper_io_base = io_base; // @[BasicChiselModules.scala 568:22]
  assign memWrapper_io_len = io_len; // @[BasicChiselModules.scala 573:21]
  assign memWrapper_io_out_ready = io_streamOut_ready; // @[BasicChiselModules.scala 575:21]
  assign memWrapper_io_start = io_start; // @[BasicChiselModules.scala 569:23]
  assign memWrapper_io_enqEn = io_enqEn; // @[BasicChiselModules.scala 571:23]
  assign memWrapper_io_deqEn = io_deqEn; // @[BasicChiselModules.scala 572:23]
  assign syncScheduleController_clock = clock;
  assign syncScheduleController_reset = reset;
  assign syncScheduleController_io_skewing = io_skewing; // @[BasicChiselModules.scala 582:37]
  assign syncScheduleController_io_input0 = {{24'd0}, io_inputs_0}; // @[BasicChiselModules.scala 579:36]
  assign syncScheduleController_io_input1 = io_inputs_1; // @[BasicChiselModules.scala 580:36]
endmodule
module ConfigController(
  input          clock,
  input          reset,
  input          io_en,
  input  [2:0]   io_II,
  output [779:0] io_outConfig
);
  reg  state; // @[BasicChiselModules.scala 64:22]
  reg [31:0] _RAND_0;
  reg [2:0] cycleReg; // @[BasicChiselModules.scala 65:21]
  reg [31:0] _RAND_1;
  reg [779:0] configRegs_0; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_2;
  reg [779:0] configRegs_1; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_3;
  reg [779:0] configRegs_2; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_4;
  reg [779:0] configRegs_3; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_5;
  reg [779:0] configRegs_4; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_6;
  reg [779:0] configRegs_5; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_7;
  reg [779:0] configRegs_6; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_8;
  reg [779:0] configRegs_7; // @[BasicChiselModules.scala 67:27]
  reg [799:0] _RAND_9;
  wire  _T_1; // @[BasicChiselModules.scala 71:14]
  wire [779:0] _GEN_1; // @[BasicChiselModules.scala 74:18]
  wire [779:0] _GEN_2; // @[BasicChiselModules.scala 74:18]
  wire [779:0] _GEN_3; // @[BasicChiselModules.scala 74:18]
  wire [779:0] _GEN_4; // @[BasicChiselModules.scala 74:18]
  wire [779:0] _GEN_5; // @[BasicChiselModules.scala 74:18]
  wire [779:0] _GEN_6; // @[BasicChiselModules.scala 74:18]
  wire [779:0] _GEN_7; // @[BasicChiselModules.scala 74:18]
  wire  _T_3; // @[BasicChiselModules.scala 80:21]
  wire [2:0] _T_5; // @[BasicChiselModules.scala 84:30]
  wire  _GEN_17; // @[BasicChiselModules.scala 80:31]
  wire [2:0] _T_7; // @[BasicChiselModules.scala 87:31]
  wire  _T_8; // @[BasicChiselModules.scala 87:21]
  wire  _GEN_28; // @[BasicChiselModules.scala 78:33]
  wire  _GEN_38; // @[BasicChiselModules.scala 77:14]
  assign _T_1 = state == 1'h0; // @[BasicChiselModules.scala 71:14]
  assign _GEN_1 = 3'h1 == cycleReg ? configRegs_1 : configRegs_0; // @[BasicChiselModules.scala 74:18]
  assign _GEN_2 = 3'h2 == cycleReg ? configRegs_2 : _GEN_1; // @[BasicChiselModules.scala 74:18]
  assign _GEN_3 = 3'h3 == cycleReg ? configRegs_3 : _GEN_2; // @[BasicChiselModules.scala 74:18]
  assign _GEN_4 = 3'h4 == cycleReg ? configRegs_4 : _GEN_3; // @[BasicChiselModules.scala 74:18]
  assign _GEN_5 = 3'h5 == cycleReg ? configRegs_5 : _GEN_4; // @[BasicChiselModules.scala 74:18]
  assign _GEN_6 = 3'h6 == cycleReg ? configRegs_6 : _GEN_5; // @[BasicChiselModules.scala 74:18]
  assign _GEN_7 = 3'h7 == cycleReg ? configRegs_7 : _GEN_6; // @[BasicChiselModules.scala 74:18]
  assign _T_3 = cycleReg == io_II; // @[BasicChiselModules.scala 80:21]
  assign _T_5 = cycleReg + 3'h1; // @[BasicChiselModules.scala 84:30]
  assign _GEN_17 = _T_3 | state; // @[BasicChiselModules.scala 80:31]
  assign _T_7 = io_II - 3'h1; // @[BasicChiselModules.scala 87:31]
  assign _T_8 = cycleReg == _T_7; // @[BasicChiselModules.scala 87:21]
  assign _GEN_28 = _T_1 ? _GEN_17 : state; // @[BasicChiselModules.scala 78:33]
  assign _GEN_38 = io_en & _GEN_28; // @[BasicChiselModules.scala 77:14]
  assign io_outConfig = _T_1 ? 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d : _GEN_7; // @[BasicChiselModules.scala 72:18 BasicChiselModules.scala 74:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cycleReg = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {25{`RANDOM}};
  configRegs_0 = _RAND_2[779:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {25{`RANDOM}};
  configRegs_1 = _RAND_3[779:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {25{`RANDOM}};
  configRegs_2 = _RAND_4[779:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {25{`RANDOM}};
  configRegs_3 = _RAND_5[779:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {25{`RANDOM}};
  configRegs_4 = _RAND_6[779:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {25{`RANDOM}};
  configRegs_5 = _RAND_7[779:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {25{`RANDOM}};
  configRegs_6 = _RAND_8[779:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {25{`RANDOM}};
  configRegs_7 = _RAND_9[779:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      state <= _GEN_38;
    end
    if (io_en) begin
      if (_T_1) begin
        if (_T_3) begin
          cycleReg <= 3'h0;
        end else begin
          cycleReg <= _T_5;
        end
      end else if (_T_8) begin
        cycleReg <= 3'h0;
      end else begin
        cycleReg <= _T_5;
      end
    end else begin
      cycleReg <= 3'h0;
    end
    if (reset) begin
      configRegs_0 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h0 == cycleReg) begin
          configRegs_0 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
    if (reset) begin
      configRegs_1 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h1 == cycleReg) begin
          configRegs_1 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
    if (reset) begin
      configRegs_2 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h2 == cycleReg) begin
          configRegs_2 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
    if (reset) begin
      configRegs_3 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h3 == cycleReg) begin
          configRegs_3 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
    if (reset) begin
      configRegs_4 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h4 == cycleReg) begin
          configRegs_4 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
    if (reset) begin
      configRegs_5 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h5 == cycleReg) begin
          configRegs_5 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
    if (reset) begin
      configRegs_6 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h6 == cycleReg) begin
          configRegs_6 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
    if (reset) begin
      configRegs_7 <= 780'h0;
    end else if (io_en) begin
      if (_T_1) begin
        if (3'h7 == cycleReg) begin
          configRegs_7 <= 780'h15940000000001a0000000008c000000000864b000080694000000003b80000000011b00000000000030000000088000000000dc0000000001a0a20000000042e80000000000007700000000081a000000000000000000bb54000000020d;
        end
      end
    end
  end
endmodule
module Dispatch_14(
  input         io_en,
  input  [41:0] io_configuration,
  output [31:0] io_outs_3,
  output [2:0]  io_outs_2,
  output [2:0]  io_outs_1,
  output [3:0]  io_outs_0
);
  wire [3:0] _T; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_1; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_2; // @[BasicChiselModules.scala 409:37]
  wire [31:0] _T_3; // @[BasicChiselModules.scala 409:37]
  assign _T = io_configuration[3:0]; // @[BasicChiselModules.scala 409:37]
  assign _T_1 = io_configuration[6:4]; // @[BasicChiselModules.scala 409:37]
  assign _T_2 = io_configuration[9:7]; // @[BasicChiselModules.scala 409:37]
  assign _T_3 = io_configuration[41:10]; // @[BasicChiselModules.scala 409:37]
  assign io_outs_3 = io_en ? _T_3 : 32'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_2 = io_en ? _T_2 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_1 = io_en ? _T_1 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_0 = io_en ? _T : 4'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module Dispatch_15(
  input         io_en,
  input  [44:0] io_configuration,
  output [31:0] io_outs_4,
  output [2:0]  io_outs_3,
  output [2:0]  io_outs_2,
  output [2:0]  io_outs_1,
  output [3:0]  io_outs_0
);
  wire [3:0] _T; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_1; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_2; // @[BasicChiselModules.scala 409:37]
  wire [2:0] _T_3; // @[BasicChiselModules.scala 409:37]
  wire [31:0] _T_4; // @[BasicChiselModules.scala 409:37]
  assign _T = io_configuration[3:0]; // @[BasicChiselModules.scala 409:37]
  assign _T_1 = io_configuration[6:4]; // @[BasicChiselModules.scala 409:37]
  assign _T_2 = io_configuration[9:7]; // @[BasicChiselModules.scala 409:37]
  assign _T_3 = io_configuration[12:10]; // @[BasicChiselModules.scala 409:37]
  assign _T_4 = io_configuration[44:13]; // @[BasicChiselModules.scala 409:37]
  assign io_outs_4 = io_en ? _T_4 : 32'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_3 = io_en ? _T_3 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_2 = io_en ? _T_2 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_1 = io_en ? _T_1 : 3'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_0 = io_en ? _T : 4'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module Dispatch_19(
  input         io_en,
  input  [15:0] io_configuration,
  output [1:0]  io_outs_7,
  output [1:0]  io_outs_6,
  output [1:0]  io_outs_5,
  output [1:0]  io_outs_4,
  output [1:0]  io_outs_3,
  output [1:0]  io_outs_2,
  output [1:0]  io_outs_1,
  output [1:0]  io_outs_0
);
  wire [1:0] _T; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_1; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_2; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_3; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_4; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_5; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_6; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_7; // @[BasicChiselModules.scala 409:37]
  assign _T = io_configuration[1:0]; // @[BasicChiselModules.scala 409:37]
  assign _T_1 = io_configuration[3:2]; // @[BasicChiselModules.scala 409:37]
  assign _T_2 = io_configuration[5:4]; // @[BasicChiselModules.scala 409:37]
  assign _T_3 = io_configuration[7:6]; // @[BasicChiselModules.scala 409:37]
  assign _T_4 = io_configuration[9:8]; // @[BasicChiselModules.scala 409:37]
  assign _T_5 = io_configuration[11:10]; // @[BasicChiselModules.scala 409:37]
  assign _T_6 = io_configuration[13:12]; // @[BasicChiselModules.scala 409:37]
  assign _T_7 = io_configuration[15:14]; // @[BasicChiselModules.scala 409:37]
  assign io_outs_7 = io_en ? _T_7 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_6 = io_en ? _T_6 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_5 = io_en ? _T_5 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_4 = io_en ? _T_4 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_3 = io_en ? _T_3 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_2 = io_en ? _T_2 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_1 = io_en ? _T_1 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_0 = io_en ? _T : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module Dispatch_21(
  input        io_en,
  input  [4:0] io_configuration,
  output       io_outs_2,
  output [1:0] io_outs_1,
  output [1:0] io_outs_0
);
  wire [1:0] _T; // @[BasicChiselModules.scala 409:37]
  wire [1:0] _T_1; // @[BasicChiselModules.scala 409:37]
  wire  _T_2; // @[BasicChiselModules.scala 409:37]
  assign _T = io_configuration[1:0]; // @[BasicChiselModules.scala 409:37]
  assign _T_1 = io_configuration[3:2]; // @[BasicChiselModules.scala 409:37]
  assign _T_2 = io_configuration[4]; // @[BasicChiselModules.scala 409:37]
  assign io_outs_2 = io_en & _T_2; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_1 = io_en ? _T_1 : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_0 = io_en ? _T : 2'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module Dispatch_30(
  input         io_en,
  input  [35:0] io_configuration,
  output [35:0] io_outs_0
);
  assign io_outs_0 = io_en ? io_configuration : 36'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module Dispatch_36(
  input          io_en,
  input  [779:0] io_configuration,
  output [41:0]  io_outs_21,
  output [44:0]  io_outs_20,
  output [44:0]  io_outs_19,
  output [44:0]  io_outs_18,
  output [4:0]   io_outs_17,
  output [35:0]  io_outs_16,
  output [44:0]  io_outs_15,
  output [4:0]   io_outs_14,
  output [41:0]  io_outs_13,
  output [44:0]  io_outs_12,
  output [4:0]   io_outs_11,
  output [44:0]  io_outs_10,
  output [44:0]  io_outs_9,
  output [44:0]  io_outs_8,
  output [4:0]   io_outs_7,
  output [44:0]  io_outs_6,
  output [15:0]  io_outs_5,
  output [44:0]  io_outs_4,
  output [44:0]  io_outs_3,
  output [41:0]  io_outs_2,
  output [44:0]  io_outs_1,
  output [41:0]  io_outs_0
);
  wire [41:0] _T; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_1; // @[BasicChiselModules.scala 409:37]
  wire [41:0] _T_2; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_3; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_4; // @[BasicChiselModules.scala 409:37]
  wire [15:0] _T_5; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_6; // @[BasicChiselModules.scala 409:37]
  wire [4:0] _T_7; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_8; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_9; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_10; // @[BasicChiselModules.scala 409:37]
  wire [4:0] _T_11; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_12; // @[BasicChiselModules.scala 409:37]
  wire [41:0] _T_13; // @[BasicChiselModules.scala 409:37]
  wire [4:0] _T_14; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_15; // @[BasicChiselModules.scala 409:37]
  wire [35:0] _T_16; // @[BasicChiselModules.scala 409:37]
  wire [4:0] _T_17; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_18; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_19; // @[BasicChiselModules.scala 409:37]
  wire [44:0] _T_20; // @[BasicChiselModules.scala 409:37]
  wire [41:0] _T_21; // @[BasicChiselModules.scala 409:37]
  assign _T = io_configuration[41:0]; // @[BasicChiselModules.scala 409:37]
  assign _T_1 = io_configuration[86:42]; // @[BasicChiselModules.scala 409:37]
  assign _T_2 = io_configuration[128:87]; // @[BasicChiselModules.scala 409:37]
  assign _T_3 = io_configuration[173:129]; // @[BasicChiselModules.scala 409:37]
  assign _T_4 = io_configuration[218:174]; // @[BasicChiselModules.scala 409:37]
  assign _T_5 = io_configuration[234:219]; // @[BasicChiselModules.scala 409:37]
  assign _T_6 = io_configuration[279:235]; // @[BasicChiselModules.scala 409:37]
  assign _T_7 = io_configuration[284:280]; // @[BasicChiselModules.scala 409:37]
  assign _T_8 = io_configuration[329:285]; // @[BasicChiselModules.scala 409:37]
  assign _T_9 = io_configuration[374:330]; // @[BasicChiselModules.scala 409:37]
  assign _T_10 = io_configuration[419:375]; // @[BasicChiselModules.scala 409:37]
  assign _T_11 = io_configuration[424:420]; // @[BasicChiselModules.scala 409:37]
  assign _T_12 = io_configuration[469:425]; // @[BasicChiselModules.scala 409:37]
  assign _T_13 = io_configuration[511:470]; // @[BasicChiselModules.scala 409:37]
  assign _T_14 = io_configuration[516:512]; // @[BasicChiselModules.scala 409:37]
  assign _T_15 = io_configuration[561:517]; // @[BasicChiselModules.scala 409:37]
  assign _T_16 = io_configuration[597:562]; // @[BasicChiselModules.scala 409:37]
  assign _T_17 = io_configuration[602:598]; // @[BasicChiselModules.scala 409:37]
  assign _T_18 = io_configuration[647:603]; // @[BasicChiselModules.scala 409:37]
  assign _T_19 = io_configuration[692:648]; // @[BasicChiselModules.scala 409:37]
  assign _T_20 = io_configuration[737:693]; // @[BasicChiselModules.scala 409:37]
  assign _T_21 = io_configuration[779:738]; // @[BasicChiselModules.scala 409:37]
  assign io_outs_21 = io_en ? _T_21 : 42'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_20 = io_en ? _T_20 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_19 = io_en ? _T_19 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_18 = io_en ? _T_18 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_17 = io_en ? _T_17 : 5'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_16 = io_en ? _T_16 : 36'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_15 = io_en ? _T_15 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_14 = io_en ? _T_14 : 5'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_13 = io_en ? _T_13 : 42'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_12 = io_en ? _T_12 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_11 = io_en ? _T_11 : 5'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_10 = io_en ? _T_10 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_9 = io_en ? _T_9 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_8 = io_en ? _T_8 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_7 = io_en ? _T_7 : 5'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_6 = io_en ? _T_6 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_5 = io_en ? _T_5 : 16'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_4 = io_en ? _T_4 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_3 = io_en ? _T_3 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_2 = io_en ? _T_2 : 42'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_1 = io_en ? _T_1 : 45'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
  assign io_outs_0 = io_en ? _T : 42'h0; // @[BasicChiselModules.scala 409:18 BasicChiselModules.scala 415:11]
endmodule
module TopModule(
  input         clock,
  input         reset,
  output        io_streamInLSU_3_ready,
  input         io_streamInLSU_3_valid,
  input  [31:0] io_streamInLSU_3_bits,
  output        io_streamInLSU_2_ready,
  input         io_streamInLSU_2_valid,
  input  [31:0] io_streamInLSU_2_bits,
  output        io_streamInLSU_1_ready,
  input         io_streamInLSU_1_valid,
  input  [31:0] io_streamInLSU_1_bits,
  output        io_streamInLSU_0_ready,
  input         io_streamInLSU_0_valid,
  input  [31:0] io_streamInLSU_0_bits,
  input         io_streamOutLSU_3_ready,
  output        io_streamOutLSU_3_valid,
  output [31:0] io_streamOutLSU_3_bits,
  input         io_streamOutLSU_2_ready,
  output        io_streamOutLSU_2_valid,
  output [31:0] io_streamOutLSU_2_bits,
  input         io_streamOutLSU_1_ready,
  output        io_streamOutLSU_1_valid,
  output [31:0] io_streamOutLSU_1_bits,
  input         io_streamOutLSU_0_ready,
  output        io_streamOutLSU_0_valid,
  output [31:0] io_streamOutLSU_0_bits,
  input  [7:0]  io_baseLSU_0,
  input  [7:0]  io_baseLSU_1,
  input  [7:0]  io_baseLSU_2,
  input  [7:0]  io_baseLSU_3,
  input  [7:0]  io_lenLSU_0,
  input  [7:0]  io_lenLSU_1,
  input  [7:0]  io_lenLSU_2,
  input  [7:0]  io_lenLSU_3,
  input         io_startLSU_0,
  input         io_startLSU_1,
  input         io_startLSU_2,
  input         io_startLSU_3,
  input         io_enqEnLSU_0,
  input         io_enqEnLSU_1,
  input         io_enqEnLSU_2,
  input         io_enqEnLSU_3,
  input         io_deqEnLSU_0,
  input         io_deqEnLSU_1,
  input         io_deqEnLSU_2,
  input         io_deqEnLSU_3,
  output        io_idleLSU_0,
  output        io_idleLSU_1,
  output        io_idleLSU_2,
  output        io_idleLSU_3,
  input         io_en,
  input  [2:0]  io_II,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_3,
  output [31:0] io_outs_2,
  output [31:0] io_outs_1,
  output [31:0] io_outs_0
);
  wire  scheduleDispatch_io_en; // @[TopModule.scala 119:32]
  wire [8:0] scheduleDispatch_io_outs_144; // @[TopModule.scala 119:32]
  wire  Alu_clock; // @[TopModule.scala 123:54]
  wire  Alu_reset; // @[TopModule.scala 123:54]
  wire  Alu_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_1_clock; // @[TopModule.scala 123:54]
  wire  Alu_1_reset; // @[TopModule.scala 123:54]
  wire  Alu_1_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_1_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_1_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_1_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_1_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_1_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_2_clock; // @[TopModule.scala 123:54]
  wire  Alu_2_reset; // @[TopModule.scala 123:54]
  wire  Alu_2_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_2_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_2_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_2_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_2_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_2_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_3_clock; // @[TopModule.scala 123:54]
  wire  Alu_3_reset; // @[TopModule.scala 123:54]
  wire  Alu_3_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_3_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_3_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_3_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_3_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_3_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_4_clock; // @[TopModule.scala 123:54]
  wire  Alu_4_reset; // @[TopModule.scala 123:54]
  wire  Alu_4_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_4_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_4_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_4_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_4_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_4_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_5_clock; // @[TopModule.scala 123:54]
  wire  Alu_5_reset; // @[TopModule.scala 123:54]
  wire  Alu_5_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_5_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_5_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_5_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_5_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_5_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_6_clock; // @[TopModule.scala 123:54]
  wire  Alu_6_reset; // @[TopModule.scala 123:54]
  wire  Alu_6_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_6_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_6_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_6_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_6_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_6_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_7_clock; // @[TopModule.scala 123:54]
  wire  Alu_7_reset; // @[TopModule.scala 123:54]
  wire  Alu_7_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_7_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_7_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_7_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_7_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_7_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_8_clock; // @[TopModule.scala 123:54]
  wire  Alu_8_reset; // @[TopModule.scala 123:54]
  wire  Alu_8_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_8_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_8_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_8_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_8_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_8_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_9_clock; // @[TopModule.scala 123:54]
  wire  Alu_9_reset; // @[TopModule.scala 123:54]
  wire  Alu_9_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_9_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_9_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_9_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_9_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_9_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_10_clock; // @[TopModule.scala 123:54]
  wire  Alu_10_reset; // @[TopModule.scala 123:54]
  wire  Alu_10_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_10_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_10_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_10_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_10_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_10_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_11_clock; // @[TopModule.scala 123:54]
  wire  Alu_11_reset; // @[TopModule.scala 123:54]
  wire  Alu_11_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_11_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_11_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_11_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_11_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_11_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_12_clock; // @[TopModule.scala 123:54]
  wire  Alu_12_reset; // @[TopModule.scala 123:54]
  wire  Alu_12_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_12_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_12_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_12_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_12_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_12_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_13_clock; // @[TopModule.scala 123:54]
  wire  Alu_13_reset; // @[TopModule.scala 123:54]
  wire  Alu_13_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_13_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_13_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_13_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_13_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_13_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_14_clock; // @[TopModule.scala 123:54]
  wire  Alu_14_reset; // @[TopModule.scala 123:54]
  wire  Alu_14_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_14_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_14_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_14_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_14_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_14_io_outs_0; // @[TopModule.scala 123:54]
  wire  Alu_15_clock; // @[TopModule.scala 123:54]
  wire  Alu_15_reset; // @[TopModule.scala 123:54]
  wire  Alu_15_io_en; // @[TopModule.scala 123:54]
  wire [4:0] Alu_15_io_skewing; // @[TopModule.scala 123:54]
  wire [3:0] Alu_15_io_configuration; // @[TopModule.scala 123:54]
  wire [31:0] Alu_15_io_inputs_1; // @[TopModule.scala 123:54]
  wire [31:0] Alu_15_io_inputs_0; // @[TopModule.scala 123:54]
  wire [31:0] Alu_15_io_outs_0; // @[TopModule.scala 123:54]
  wire  MultiIIScheduleController_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_1_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_1_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_1_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_1_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_1_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_1_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_2_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_2_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_2_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_2_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_2_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_2_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_3_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_3_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_3_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_3_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_3_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_3_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_4_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_4_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_4_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_4_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_4_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_4_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_4_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_5_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_5_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_5_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_5_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_5_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_5_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_5_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_6_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_6_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_6_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_6_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_6_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_6_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_6_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_7_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_7_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_7_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_7_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_7_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_7_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_7_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_8_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_8_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_8_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_8_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_8_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_8_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_8_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_9_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_9_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_9_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_9_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_9_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_9_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_9_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_10_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_10_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_10_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_10_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_10_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_10_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_10_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_11_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_11_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_11_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_11_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_11_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_11_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_11_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_12_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_12_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_12_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_12_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_12_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_12_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_12_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_13_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_13_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_13_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_13_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_13_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_13_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_13_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_14_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_14_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_14_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_14_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_14_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_14_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_14_io_skewing; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_15_clock; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_15_reset; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_15_io_en; // @[TopModule.scala 125:72]
  wire [8:0] MultiIIScheduleController_15_io_schedules_0; // @[TopModule.scala 125:72]
  wire [2:0] MultiIIScheduleController_15_io_II; // @[TopModule.scala 125:72]
  wire  MultiIIScheduleController_15_io_valid; // @[TopModule.scala 125:72]
  wire [4:0] MultiIIScheduleController_15_io_skewing; // @[TopModule.scala 125:72]
  wire  RegisterFiles_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_io_en; // @[TopModule.scala 143:21]
  wire [35:0] RegisterFiles_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_inputs_3; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_inputs_2; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_inputs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_7; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_6; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_5; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_4; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_3; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_2; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_1_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_1_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_1_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_1_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_1_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_1_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_1_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_2_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_2_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_2_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_2_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_2_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_2_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_2_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_3_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_3_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_3_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_3_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_3_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_3_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_3_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_4_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_4_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_4_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_4_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_4_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_4_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_4_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_5_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_5_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_5_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_5_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_5_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_5_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_5_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_6_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_6_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_6_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_6_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_6_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_6_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_6_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_7_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_7_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_7_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_7_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_7_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_7_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_7_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_8_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_8_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_8_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_8_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_8_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_8_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_8_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_9_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_9_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_9_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_9_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_9_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_9_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_9_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_10_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_10_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_10_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_10_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_10_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_10_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_10_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_11_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_11_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_11_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_11_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_11_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_11_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_11_io_outs_0; // @[TopModule.scala 143:21]
  wire  RegisterFiles_12_clock; // @[TopModule.scala 143:21]
  wire  RegisterFiles_12_reset; // @[TopModule.scala 143:21]
  wire  RegisterFiles_12_io_en; // @[TopModule.scala 143:21]
  wire [2:0] RegisterFiles_12_io_configuration; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_12_io_inputs_0; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_12_io_outs_1; // @[TopModule.scala 143:21]
  wire [31:0] RegisterFiles_12_io_outs_0; // @[TopModule.scala 143:21]
  wire  Multiplexer_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_1_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_1_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_1_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_1_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_1_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_1_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_1_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_2_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_2_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_2_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_2_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_2_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_2_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_2_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_3_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_3_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_3_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_3_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_3_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_3_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_3_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_4_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_4_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_4_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_4_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_4_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_4_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_4_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_5_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_5_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_5_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_5_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_5_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_5_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_5_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_6_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_6_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_6_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_6_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_6_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_6_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_6_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_7_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_7_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_7_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_7_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_7_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_7_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_7_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_8_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_8_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_7; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_8_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_9_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_9_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_9_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_10_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_10_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_7; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_10_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_11_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_11_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_11_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_12_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_12_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_7; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_12_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_13_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_13_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_13_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_14_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_14_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_7; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_14_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_15_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_15_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_15_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_16_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_16_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_16_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_17_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_17_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_17_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_17_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_17_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_17_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_17_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_17_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_17_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_18_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_18_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_18_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_19_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_19_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_19_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_19_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_19_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_19_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_19_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_19_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_19_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_20_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_20_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_20_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_21_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_21_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_21_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_21_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_21_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_21_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_21_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_21_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_21_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_22_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_22_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_22_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_23_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_23_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_23_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_23_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_23_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_23_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_23_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_23_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_23_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_24_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_24_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_24_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_25_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_25_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_25_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_25_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_25_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_25_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_25_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_25_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_25_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_26_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_26_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_26_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_27_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_27_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_27_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_27_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_27_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_27_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_27_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_27_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_27_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_28_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_28_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_28_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_29_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_29_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_29_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_29_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_29_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_29_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_29_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_29_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_29_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_30_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_30_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_30_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_31_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_31_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_31_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_31_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_31_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_31_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_31_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_31_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_31_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_32_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_32_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_32_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_33_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_33_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_33_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_33_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_33_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_33_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_33_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_33_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_33_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_34_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_34_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_34_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_35_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_35_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_35_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_35_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_35_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_35_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_35_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_35_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_35_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_36_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_36_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_36_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_37_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_37_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_37_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_37_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_37_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_37_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_37_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_37_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_37_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_38_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_38_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_inputs_6; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_38_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_39_io_en; // @[TopModule.scala 154:11]
  wire [2:0] Multiplexer_39_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_39_io_inputs_5; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_39_io_inputs_4; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_39_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_39_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_39_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_39_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_39_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_40_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_40_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_40_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_40_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_40_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_40_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_40_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_41_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_41_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_41_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_41_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_41_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_41_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_41_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_42_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_42_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_42_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_42_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_42_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_42_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_42_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_43_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_43_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_43_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_43_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_43_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_43_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_43_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_44_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_44_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_44_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_44_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_44_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_44_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_44_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_45_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_45_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_45_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_45_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_45_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_45_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_45_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_46_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_46_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_46_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_46_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_46_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_46_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_46_io_outs_0; // @[TopModule.scala 154:11]
  wire  Multiplexer_47_io_en; // @[TopModule.scala 154:11]
  wire [1:0] Multiplexer_47_io_configuration; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_47_io_inputs_3; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_47_io_inputs_2; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_47_io_inputs_1; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_47_io_inputs_0; // @[TopModule.scala 154:11]
  wire [31:0] Multiplexer_47_io_outs_0; // @[TopModule.scala 154:11]
  wire  ConstUnit_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_1_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_1_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_1_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_2_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_2_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_2_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_3_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_3_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_3_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_4_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_4_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_4_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_5_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_5_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_5_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_6_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_6_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_6_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_7_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_7_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_7_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_8_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_8_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_8_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_9_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_9_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_9_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_10_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_10_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_10_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_11_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_11_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_11_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_12_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_12_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_12_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_13_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_13_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_13_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_14_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_14_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_14_io_outs_0; // @[TopModule.scala 163:21]
  wire  ConstUnit_15_io_en; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_15_io_configuration; // @[TopModule.scala 163:21]
  wire [31:0] ConstUnit_15_io_outs_0; // @[TopModule.scala 163:21]
  wire  LoadStoreUnit_clock; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_reset; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_configuration; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_en; // @[TopModule.scala 171:21]
  wire [4:0] LoadStoreUnit_io_skewing; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_streamIn_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_streamIn_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_io_streamIn_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_io_len; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_streamOut_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_streamOut_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_io_streamOut_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_io_base; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_start; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_enqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_deqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_io_idle; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_io_inputs_1; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_io_inputs_0; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_io_outs_0; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_clock; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_reset; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_configuration; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_en; // @[TopModule.scala 171:21]
  wire [4:0] LoadStoreUnit_1_io_skewing; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_streamIn_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_streamIn_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_1_io_streamIn_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_1_io_len; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_streamOut_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_streamOut_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_1_io_streamOut_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_1_io_base; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_start; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_enqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_deqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_1_io_idle; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_1_io_inputs_1; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_1_io_inputs_0; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_clock; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_reset; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_configuration; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_en; // @[TopModule.scala 171:21]
  wire [4:0] LoadStoreUnit_2_io_skewing; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_streamIn_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_streamIn_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_2_io_streamIn_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_2_io_len; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_streamOut_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_streamOut_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_2_io_streamOut_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_2_io_base; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_start; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_enqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_deqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_2_io_idle; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_2_io_inputs_1; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_2_io_inputs_0; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_clock; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_reset; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_configuration; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_en; // @[TopModule.scala 171:21]
  wire [4:0] LoadStoreUnit_3_io_skewing; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_streamIn_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_streamIn_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_3_io_streamIn_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_3_io_len; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_streamOut_ready; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_streamOut_valid; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_3_io_streamOut_bits; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_3_io_base; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_start; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_enqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_deqEn; // @[TopModule.scala 171:21]
  wire  LoadStoreUnit_3_io_idle; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_3_io_inputs_1; // @[TopModule.scala 171:21]
  wire [7:0] LoadStoreUnit_3_io_inputs_0; // @[TopModule.scala 171:21]
  wire [31:0] LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 171:21]
  wire  MultiIIScheduleController_16_clock; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_16_reset; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_16_io_en; // @[TopModule.scala 172:78]
  wire [8:0] MultiIIScheduleController_16_io_schedules_0; // @[TopModule.scala 172:78]
  wire [2:0] MultiIIScheduleController_16_io_II; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_16_io_valid; // @[TopModule.scala 172:78]
  wire [4:0] MultiIIScheduleController_16_io_skewing; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_17_clock; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_17_reset; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_17_io_en; // @[TopModule.scala 172:78]
  wire [8:0] MultiIIScheduleController_17_io_schedules_0; // @[TopModule.scala 172:78]
  wire [2:0] MultiIIScheduleController_17_io_II; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_17_io_valid; // @[TopModule.scala 172:78]
  wire [4:0] MultiIIScheduleController_17_io_skewing; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_18_clock; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_18_reset; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_18_io_en; // @[TopModule.scala 172:78]
  wire [8:0] MultiIIScheduleController_18_io_schedules_0; // @[TopModule.scala 172:78]
  wire [2:0] MultiIIScheduleController_18_io_II; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_18_io_valid; // @[TopModule.scala 172:78]
  wire [4:0] MultiIIScheduleController_18_io_skewing; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_19_clock; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_19_reset; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_19_io_en; // @[TopModule.scala 172:78]
  wire [8:0] MultiIIScheduleController_19_io_schedules_0; // @[TopModule.scala 172:78]
  wire [2:0] MultiIIScheduleController_19_io_II; // @[TopModule.scala 172:78]
  wire  MultiIIScheduleController_19_io_valid; // @[TopModule.scala 172:78]
  wire [4:0] MultiIIScheduleController_19_io_skewing; // @[TopModule.scala 172:78]
  wire  configController_clock; // @[TopModule.scala 219:32]
  wire  configController_reset; // @[TopModule.scala 219:32]
  wire  configController_io_en; // @[TopModule.scala 219:32]
  wire [2:0] configController_io_II; // @[TopModule.scala 219:32]
  wire [779:0] configController_io_outConfig; // @[TopModule.scala 219:32]
  wire  dispatchs_0_io_en; // @[TopModule.scala 246:26]
  wire [41:0] dispatchs_0_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_0_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_0_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_0_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_0_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_1_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_1_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_1_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_1_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_1_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_1_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_1_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_2_io_en; // @[TopModule.scala 246:26]
  wire [41:0] dispatchs_2_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_2_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_2_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_2_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_2_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_3_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_3_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_3_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_3_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_3_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_3_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_3_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_4_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_4_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_4_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_4_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_4_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_4_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_4_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_5_io_en; // @[TopModule.scala 246:26]
  wire [15:0] dispatchs_5_io_configuration; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_7; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_6; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_5; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_4; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_3; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_2; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_1; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_5_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_6_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_6_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_6_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_6_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_6_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_6_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_6_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_7_io_en; // @[TopModule.scala 246:26]
  wire [4:0] dispatchs_7_io_configuration; // @[TopModule.scala 246:26]
  wire  dispatchs_7_io_outs_2; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_7_io_outs_1; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_7_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_8_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_8_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_8_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_8_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_8_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_8_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_8_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_9_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_9_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_9_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_9_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_9_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_9_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_9_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_10_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_10_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_10_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_10_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_10_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_10_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_10_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_11_io_en; // @[TopModule.scala 246:26]
  wire [4:0] dispatchs_11_io_configuration; // @[TopModule.scala 246:26]
  wire  dispatchs_11_io_outs_2; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_11_io_outs_1; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_11_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_12_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_12_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_12_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_12_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_12_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_12_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_12_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_13_io_en; // @[TopModule.scala 246:26]
  wire [41:0] dispatchs_13_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_13_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_13_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_13_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_13_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_14_io_en; // @[TopModule.scala 246:26]
  wire [4:0] dispatchs_14_io_configuration; // @[TopModule.scala 246:26]
  wire  dispatchs_14_io_outs_2; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_14_io_outs_1; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_14_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_15_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_15_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_15_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_15_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_15_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_15_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_15_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_16_io_en; // @[TopModule.scala 246:26]
  wire [35:0] dispatchs_16_io_configuration; // @[TopModule.scala 246:26]
  wire [35:0] dispatchs_16_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_17_io_en; // @[TopModule.scala 246:26]
  wire [4:0] dispatchs_17_io_configuration; // @[TopModule.scala 246:26]
  wire  dispatchs_17_io_outs_2; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_17_io_outs_1; // @[TopModule.scala 246:26]
  wire [1:0] dispatchs_17_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_18_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_18_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_18_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_18_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_18_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_18_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_18_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_19_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_19_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_19_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_19_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_19_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_19_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_19_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_20_io_en; // @[TopModule.scala 246:26]
  wire [44:0] dispatchs_20_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_20_io_outs_4; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_20_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_20_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_20_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_20_io_outs_0; // @[TopModule.scala 246:26]
  wire  dispatchs_21_io_en; // @[TopModule.scala 246:26]
  wire [41:0] dispatchs_21_io_configuration; // @[TopModule.scala 246:26]
  wire [31:0] dispatchs_21_io_outs_3; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_21_io_outs_2; // @[TopModule.scala 246:26]
  wire [2:0] dispatchs_21_io_outs_1; // @[TopModule.scala 246:26]
  wire [3:0] dispatchs_21_io_outs_0; // @[TopModule.scala 246:26]
  wire  topDispatch_io_en; // @[TopModule.scala 255:27]
  wire [779:0] topDispatch_io_configuration; // @[TopModule.scala 255:27]
  wire [41:0] topDispatch_io_outs_21; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_20; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_19; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_18; // @[TopModule.scala 255:27]
  wire [4:0] topDispatch_io_outs_17; // @[TopModule.scala 255:27]
  wire [35:0] topDispatch_io_outs_16; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_15; // @[TopModule.scala 255:27]
  wire [4:0] topDispatch_io_outs_14; // @[TopModule.scala 255:27]
  wire [41:0] topDispatch_io_outs_13; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_12; // @[TopModule.scala 255:27]
  wire [4:0] topDispatch_io_outs_11; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_10; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_9; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_8; // @[TopModule.scala 255:27]
  wire [4:0] topDispatch_io_outs_7; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_6; // @[TopModule.scala 255:27]
  wire [15:0] topDispatch_io_outs_5; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_4; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_3; // @[TopModule.scala 255:27]
  wire [41:0] topDispatch_io_outs_2; // @[TopModule.scala 255:27]
  wire [44:0] topDispatch_io_outs_1; // @[TopModule.scala 255:27]
  wire [41:0] topDispatch_io_outs_0; // @[TopModule.scala 255:27]
  Dispatch scheduleDispatch ( // @[TopModule.scala 119:32]
    .io_en(scheduleDispatch_io_en),
    .io_outs_144(scheduleDispatch_io_outs_144)
  );
  Alu Alu ( // @[TopModule.scala 123:54]
    .clock(Alu_clock),
    .reset(Alu_reset),
    .io_en(Alu_io_en),
    .io_skewing(Alu_io_skewing),
    .io_configuration(Alu_io_configuration),
    .io_inputs_1(Alu_io_inputs_1),
    .io_inputs_0(Alu_io_inputs_0),
    .io_outs_0(Alu_io_outs_0)
  );
  Alu Alu_1 ( // @[TopModule.scala 123:54]
    .clock(Alu_1_clock),
    .reset(Alu_1_reset),
    .io_en(Alu_1_io_en),
    .io_skewing(Alu_1_io_skewing),
    .io_configuration(Alu_1_io_configuration),
    .io_inputs_1(Alu_1_io_inputs_1),
    .io_inputs_0(Alu_1_io_inputs_0),
    .io_outs_0(Alu_1_io_outs_0)
  );
  Alu Alu_2 ( // @[TopModule.scala 123:54]
    .clock(Alu_2_clock),
    .reset(Alu_2_reset),
    .io_en(Alu_2_io_en),
    .io_skewing(Alu_2_io_skewing),
    .io_configuration(Alu_2_io_configuration),
    .io_inputs_1(Alu_2_io_inputs_1),
    .io_inputs_0(Alu_2_io_inputs_0),
    .io_outs_0(Alu_2_io_outs_0)
  );
  Alu Alu_3 ( // @[TopModule.scala 123:54]
    .clock(Alu_3_clock),
    .reset(Alu_3_reset),
    .io_en(Alu_3_io_en),
    .io_skewing(Alu_3_io_skewing),
    .io_configuration(Alu_3_io_configuration),
    .io_inputs_1(Alu_3_io_inputs_1),
    .io_inputs_0(Alu_3_io_inputs_0),
    .io_outs_0(Alu_3_io_outs_0)
  );
  Alu_4 Alu_4 ( // @[TopModule.scala 123:54]
    .clock(Alu_4_clock),
    .reset(Alu_4_reset),
    .io_en(Alu_4_io_en),
    .io_skewing(Alu_4_io_skewing),
    .io_configuration(Alu_4_io_configuration),
    .io_inputs_1(Alu_4_io_inputs_1),
    .io_inputs_0(Alu_4_io_inputs_0),
    .io_outs_0(Alu_4_io_outs_0)
  );
  Alu_4 Alu_5 ( // @[TopModule.scala 123:54]
    .clock(Alu_5_clock),
    .reset(Alu_5_reset),
    .io_en(Alu_5_io_en),
    .io_skewing(Alu_5_io_skewing),
    .io_configuration(Alu_5_io_configuration),
    .io_inputs_1(Alu_5_io_inputs_1),
    .io_inputs_0(Alu_5_io_inputs_0),
    .io_outs_0(Alu_5_io_outs_0)
  );
  Alu_4 Alu_6 ( // @[TopModule.scala 123:54]
    .clock(Alu_6_clock),
    .reset(Alu_6_reset),
    .io_en(Alu_6_io_en),
    .io_skewing(Alu_6_io_skewing),
    .io_configuration(Alu_6_io_configuration),
    .io_inputs_1(Alu_6_io_inputs_1),
    .io_inputs_0(Alu_6_io_inputs_0),
    .io_outs_0(Alu_6_io_outs_0)
  );
  Alu_4 Alu_7 ( // @[TopModule.scala 123:54]
    .clock(Alu_7_clock),
    .reset(Alu_7_reset),
    .io_en(Alu_7_io_en),
    .io_skewing(Alu_7_io_skewing),
    .io_configuration(Alu_7_io_configuration),
    .io_inputs_1(Alu_7_io_inputs_1),
    .io_inputs_0(Alu_7_io_inputs_0),
    .io_outs_0(Alu_7_io_outs_0)
  );
  Alu_4 Alu_8 ( // @[TopModule.scala 123:54]
    .clock(Alu_8_clock),
    .reset(Alu_8_reset),
    .io_en(Alu_8_io_en),
    .io_skewing(Alu_8_io_skewing),
    .io_configuration(Alu_8_io_configuration),
    .io_inputs_1(Alu_8_io_inputs_1),
    .io_inputs_0(Alu_8_io_inputs_0),
    .io_outs_0(Alu_8_io_outs_0)
  );
  Alu_4 Alu_9 ( // @[TopModule.scala 123:54]
    .clock(Alu_9_clock),
    .reset(Alu_9_reset),
    .io_en(Alu_9_io_en),
    .io_skewing(Alu_9_io_skewing),
    .io_configuration(Alu_9_io_configuration),
    .io_inputs_1(Alu_9_io_inputs_1),
    .io_inputs_0(Alu_9_io_inputs_0),
    .io_outs_0(Alu_9_io_outs_0)
  );
  Alu_4 Alu_10 ( // @[TopModule.scala 123:54]
    .clock(Alu_10_clock),
    .reset(Alu_10_reset),
    .io_en(Alu_10_io_en),
    .io_skewing(Alu_10_io_skewing),
    .io_configuration(Alu_10_io_configuration),
    .io_inputs_1(Alu_10_io_inputs_1),
    .io_inputs_0(Alu_10_io_inputs_0),
    .io_outs_0(Alu_10_io_outs_0)
  );
  Alu_4 Alu_11 ( // @[TopModule.scala 123:54]
    .clock(Alu_11_clock),
    .reset(Alu_11_reset),
    .io_en(Alu_11_io_en),
    .io_skewing(Alu_11_io_skewing),
    .io_configuration(Alu_11_io_configuration),
    .io_inputs_1(Alu_11_io_inputs_1),
    .io_inputs_0(Alu_11_io_inputs_0),
    .io_outs_0(Alu_11_io_outs_0)
  );
  Alu_4 Alu_12 ( // @[TopModule.scala 123:54]
    .clock(Alu_12_clock),
    .reset(Alu_12_reset),
    .io_en(Alu_12_io_en),
    .io_skewing(Alu_12_io_skewing),
    .io_configuration(Alu_12_io_configuration),
    .io_inputs_1(Alu_12_io_inputs_1),
    .io_inputs_0(Alu_12_io_inputs_0),
    .io_outs_0(Alu_12_io_outs_0)
  );
  Alu_4 Alu_13 ( // @[TopModule.scala 123:54]
    .clock(Alu_13_clock),
    .reset(Alu_13_reset),
    .io_en(Alu_13_io_en),
    .io_skewing(Alu_13_io_skewing),
    .io_configuration(Alu_13_io_configuration),
    .io_inputs_1(Alu_13_io_inputs_1),
    .io_inputs_0(Alu_13_io_inputs_0),
    .io_outs_0(Alu_13_io_outs_0)
  );
  Alu_4 Alu_14 ( // @[TopModule.scala 123:54]
    .clock(Alu_14_clock),
    .reset(Alu_14_reset),
    .io_en(Alu_14_io_en),
    .io_skewing(Alu_14_io_skewing),
    .io_configuration(Alu_14_io_configuration),
    .io_inputs_1(Alu_14_io_inputs_1),
    .io_inputs_0(Alu_14_io_inputs_0),
    .io_outs_0(Alu_14_io_outs_0)
  );
  Alu_4 Alu_15 ( // @[TopModule.scala 123:54]
    .clock(Alu_15_clock),
    .reset(Alu_15_reset),
    .io_en(Alu_15_io_en),
    .io_skewing(Alu_15_io_skewing),
    .io_configuration(Alu_15_io_configuration),
    .io_inputs_1(Alu_15_io_inputs_1),
    .io_inputs_0(Alu_15_io_inputs_0),
    .io_outs_0(Alu_15_io_outs_0)
  );
  MultiIIScheduleController MultiIIScheduleController ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_clock),
    .reset(MultiIIScheduleController_reset),
    .io_en(MultiIIScheduleController_io_en),
    .io_schedules_0(MultiIIScheduleController_io_schedules_0),
    .io_II(MultiIIScheduleController_io_II),
    .io_valid(MultiIIScheduleController_io_valid),
    .io_skewing(MultiIIScheduleController_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_1 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_1_clock),
    .reset(MultiIIScheduleController_1_reset),
    .io_en(MultiIIScheduleController_1_io_en),
    .io_schedules_0(MultiIIScheduleController_1_io_schedules_0),
    .io_II(MultiIIScheduleController_1_io_II),
    .io_valid(MultiIIScheduleController_1_io_valid),
    .io_skewing(MultiIIScheduleController_1_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_2 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_2_clock),
    .reset(MultiIIScheduleController_2_reset),
    .io_en(MultiIIScheduleController_2_io_en),
    .io_schedules_0(MultiIIScheduleController_2_io_schedules_0),
    .io_II(MultiIIScheduleController_2_io_II),
    .io_valid(MultiIIScheduleController_2_io_valid),
    .io_skewing(MultiIIScheduleController_2_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_3 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_3_clock),
    .reset(MultiIIScheduleController_3_reset),
    .io_en(MultiIIScheduleController_3_io_en),
    .io_schedules_0(MultiIIScheduleController_3_io_schedules_0),
    .io_II(MultiIIScheduleController_3_io_II),
    .io_valid(MultiIIScheduleController_3_io_valid),
    .io_skewing(MultiIIScheduleController_3_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_4 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_4_clock),
    .reset(MultiIIScheduleController_4_reset),
    .io_en(MultiIIScheduleController_4_io_en),
    .io_schedules_0(MultiIIScheduleController_4_io_schedules_0),
    .io_II(MultiIIScheduleController_4_io_II),
    .io_valid(MultiIIScheduleController_4_io_valid),
    .io_skewing(MultiIIScheduleController_4_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_5 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_5_clock),
    .reset(MultiIIScheduleController_5_reset),
    .io_en(MultiIIScheduleController_5_io_en),
    .io_schedules_0(MultiIIScheduleController_5_io_schedules_0),
    .io_II(MultiIIScheduleController_5_io_II),
    .io_valid(MultiIIScheduleController_5_io_valid),
    .io_skewing(MultiIIScheduleController_5_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_6 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_6_clock),
    .reset(MultiIIScheduleController_6_reset),
    .io_en(MultiIIScheduleController_6_io_en),
    .io_schedules_0(MultiIIScheduleController_6_io_schedules_0),
    .io_II(MultiIIScheduleController_6_io_II),
    .io_valid(MultiIIScheduleController_6_io_valid),
    .io_skewing(MultiIIScheduleController_6_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_7 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_7_clock),
    .reset(MultiIIScheduleController_7_reset),
    .io_en(MultiIIScheduleController_7_io_en),
    .io_schedules_0(MultiIIScheduleController_7_io_schedules_0),
    .io_II(MultiIIScheduleController_7_io_II),
    .io_valid(MultiIIScheduleController_7_io_valid),
    .io_skewing(MultiIIScheduleController_7_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_8 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_8_clock),
    .reset(MultiIIScheduleController_8_reset),
    .io_en(MultiIIScheduleController_8_io_en),
    .io_schedules_0(MultiIIScheduleController_8_io_schedules_0),
    .io_II(MultiIIScheduleController_8_io_II),
    .io_valid(MultiIIScheduleController_8_io_valid),
    .io_skewing(MultiIIScheduleController_8_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_9 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_9_clock),
    .reset(MultiIIScheduleController_9_reset),
    .io_en(MultiIIScheduleController_9_io_en),
    .io_schedules_0(MultiIIScheduleController_9_io_schedules_0),
    .io_II(MultiIIScheduleController_9_io_II),
    .io_valid(MultiIIScheduleController_9_io_valid),
    .io_skewing(MultiIIScheduleController_9_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_10 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_10_clock),
    .reset(MultiIIScheduleController_10_reset),
    .io_en(MultiIIScheduleController_10_io_en),
    .io_schedules_0(MultiIIScheduleController_10_io_schedules_0),
    .io_II(MultiIIScheduleController_10_io_II),
    .io_valid(MultiIIScheduleController_10_io_valid),
    .io_skewing(MultiIIScheduleController_10_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_11 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_11_clock),
    .reset(MultiIIScheduleController_11_reset),
    .io_en(MultiIIScheduleController_11_io_en),
    .io_schedules_0(MultiIIScheduleController_11_io_schedules_0),
    .io_II(MultiIIScheduleController_11_io_II),
    .io_valid(MultiIIScheduleController_11_io_valid),
    .io_skewing(MultiIIScheduleController_11_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_12 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_12_clock),
    .reset(MultiIIScheduleController_12_reset),
    .io_en(MultiIIScheduleController_12_io_en),
    .io_schedules_0(MultiIIScheduleController_12_io_schedules_0),
    .io_II(MultiIIScheduleController_12_io_II),
    .io_valid(MultiIIScheduleController_12_io_valid),
    .io_skewing(MultiIIScheduleController_12_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_13 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_13_clock),
    .reset(MultiIIScheduleController_13_reset),
    .io_en(MultiIIScheduleController_13_io_en),
    .io_schedules_0(MultiIIScheduleController_13_io_schedules_0),
    .io_II(MultiIIScheduleController_13_io_II),
    .io_valid(MultiIIScheduleController_13_io_valid),
    .io_skewing(MultiIIScheduleController_13_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_14 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_14_clock),
    .reset(MultiIIScheduleController_14_reset),
    .io_en(MultiIIScheduleController_14_io_en),
    .io_schedules_0(MultiIIScheduleController_14_io_schedules_0),
    .io_II(MultiIIScheduleController_14_io_II),
    .io_valid(MultiIIScheduleController_14_io_valid),
    .io_skewing(MultiIIScheduleController_14_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_15 ( // @[TopModule.scala 125:72]
    .clock(MultiIIScheduleController_15_clock),
    .reset(MultiIIScheduleController_15_reset),
    .io_en(MultiIIScheduleController_15_io_en),
    .io_schedules_0(MultiIIScheduleController_15_io_schedules_0),
    .io_II(MultiIIScheduleController_15_io_II),
    .io_valid(MultiIIScheduleController_15_io_valid),
    .io_skewing(MultiIIScheduleController_15_io_skewing)
  );
  RegisterFiles RegisterFiles ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_clock),
    .reset(RegisterFiles_reset),
    .io_en(RegisterFiles_io_en),
    .io_configuration(RegisterFiles_io_configuration),
    .io_inputs_3(RegisterFiles_io_inputs_3),
    .io_inputs_2(RegisterFiles_io_inputs_2),
    .io_inputs_1(RegisterFiles_io_inputs_1),
    .io_inputs_0(RegisterFiles_io_inputs_0),
    .io_outs_7(RegisterFiles_io_outs_7),
    .io_outs_6(RegisterFiles_io_outs_6),
    .io_outs_5(RegisterFiles_io_outs_5),
    .io_outs_4(RegisterFiles_io_outs_4),
    .io_outs_3(RegisterFiles_io_outs_3),
    .io_outs_2(RegisterFiles_io_outs_2),
    .io_outs_1(RegisterFiles_io_outs_1),
    .io_outs_0(RegisterFiles_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_1 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_1_clock),
    .reset(RegisterFiles_1_reset),
    .io_en(RegisterFiles_1_io_en),
    .io_configuration(RegisterFiles_1_io_configuration),
    .io_inputs_0(RegisterFiles_1_io_inputs_0),
    .io_outs_1(RegisterFiles_1_io_outs_1),
    .io_outs_0(RegisterFiles_1_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_2 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_2_clock),
    .reset(RegisterFiles_2_reset),
    .io_en(RegisterFiles_2_io_en),
    .io_configuration(RegisterFiles_2_io_configuration),
    .io_inputs_0(RegisterFiles_2_io_inputs_0),
    .io_outs_1(RegisterFiles_2_io_outs_1),
    .io_outs_0(RegisterFiles_2_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_3 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_3_clock),
    .reset(RegisterFiles_3_reset),
    .io_en(RegisterFiles_3_io_en),
    .io_configuration(RegisterFiles_3_io_configuration),
    .io_inputs_0(RegisterFiles_3_io_inputs_0),
    .io_outs_1(RegisterFiles_3_io_outs_1),
    .io_outs_0(RegisterFiles_3_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_4 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_4_clock),
    .reset(RegisterFiles_4_reset),
    .io_en(RegisterFiles_4_io_en),
    .io_configuration(RegisterFiles_4_io_configuration),
    .io_inputs_0(RegisterFiles_4_io_inputs_0),
    .io_outs_1(RegisterFiles_4_io_outs_1),
    .io_outs_0(RegisterFiles_4_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_5 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_5_clock),
    .reset(RegisterFiles_5_reset),
    .io_en(RegisterFiles_5_io_en),
    .io_configuration(RegisterFiles_5_io_configuration),
    .io_inputs_0(RegisterFiles_5_io_inputs_0),
    .io_outs_1(RegisterFiles_5_io_outs_1),
    .io_outs_0(RegisterFiles_5_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_6 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_6_clock),
    .reset(RegisterFiles_6_reset),
    .io_en(RegisterFiles_6_io_en),
    .io_configuration(RegisterFiles_6_io_configuration),
    .io_inputs_0(RegisterFiles_6_io_inputs_0),
    .io_outs_1(RegisterFiles_6_io_outs_1),
    .io_outs_0(RegisterFiles_6_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_7 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_7_clock),
    .reset(RegisterFiles_7_reset),
    .io_en(RegisterFiles_7_io_en),
    .io_configuration(RegisterFiles_7_io_configuration),
    .io_inputs_0(RegisterFiles_7_io_inputs_0),
    .io_outs_1(RegisterFiles_7_io_outs_1),
    .io_outs_0(RegisterFiles_7_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_8 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_8_clock),
    .reset(RegisterFiles_8_reset),
    .io_en(RegisterFiles_8_io_en),
    .io_configuration(RegisterFiles_8_io_configuration),
    .io_inputs_0(RegisterFiles_8_io_inputs_0),
    .io_outs_1(RegisterFiles_8_io_outs_1),
    .io_outs_0(RegisterFiles_8_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_9 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_9_clock),
    .reset(RegisterFiles_9_reset),
    .io_en(RegisterFiles_9_io_en),
    .io_configuration(RegisterFiles_9_io_configuration),
    .io_inputs_0(RegisterFiles_9_io_inputs_0),
    .io_outs_1(RegisterFiles_9_io_outs_1),
    .io_outs_0(RegisterFiles_9_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_10 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_10_clock),
    .reset(RegisterFiles_10_reset),
    .io_en(RegisterFiles_10_io_en),
    .io_configuration(RegisterFiles_10_io_configuration),
    .io_inputs_0(RegisterFiles_10_io_inputs_0),
    .io_outs_1(RegisterFiles_10_io_outs_1),
    .io_outs_0(RegisterFiles_10_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_11 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_11_clock),
    .reset(RegisterFiles_11_reset),
    .io_en(RegisterFiles_11_io_en),
    .io_configuration(RegisterFiles_11_io_configuration),
    .io_inputs_0(RegisterFiles_11_io_inputs_0),
    .io_outs_1(RegisterFiles_11_io_outs_1),
    .io_outs_0(RegisterFiles_11_io_outs_0)
  );
  RegisterFiles_1 RegisterFiles_12 ( // @[TopModule.scala 143:21]
    .clock(RegisterFiles_12_clock),
    .reset(RegisterFiles_12_reset),
    .io_en(RegisterFiles_12_io_en),
    .io_configuration(RegisterFiles_12_io_configuration),
    .io_inputs_0(RegisterFiles_12_io_inputs_0),
    .io_outs_1(RegisterFiles_12_io_outs_1),
    .io_outs_0(RegisterFiles_12_io_outs_0)
  );
  Multiplexer Multiplexer ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_io_en),
    .io_configuration(Multiplexer_io_configuration),
    .io_inputs_3(Multiplexer_io_inputs_3),
    .io_inputs_2(Multiplexer_io_inputs_2),
    .io_inputs_1(Multiplexer_io_inputs_1),
    .io_inputs_0(Multiplexer_io_inputs_0),
    .io_outs_0(Multiplexer_io_outs_0)
  );
  Multiplexer Multiplexer_1 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_1_io_en),
    .io_configuration(Multiplexer_1_io_configuration),
    .io_inputs_3(Multiplexer_1_io_inputs_3),
    .io_inputs_2(Multiplexer_1_io_inputs_2),
    .io_inputs_1(Multiplexer_1_io_inputs_1),
    .io_inputs_0(Multiplexer_1_io_inputs_0),
    .io_outs_0(Multiplexer_1_io_outs_0)
  );
  Multiplexer Multiplexer_2 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_2_io_en),
    .io_configuration(Multiplexer_2_io_configuration),
    .io_inputs_3(Multiplexer_2_io_inputs_3),
    .io_inputs_2(Multiplexer_2_io_inputs_2),
    .io_inputs_1(Multiplexer_2_io_inputs_1),
    .io_inputs_0(Multiplexer_2_io_inputs_0),
    .io_outs_0(Multiplexer_2_io_outs_0)
  );
  Multiplexer Multiplexer_3 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_3_io_en),
    .io_configuration(Multiplexer_3_io_configuration),
    .io_inputs_3(Multiplexer_3_io_inputs_3),
    .io_inputs_2(Multiplexer_3_io_inputs_2),
    .io_inputs_1(Multiplexer_3_io_inputs_1),
    .io_inputs_0(Multiplexer_3_io_inputs_0),
    .io_outs_0(Multiplexer_3_io_outs_0)
  );
  Multiplexer Multiplexer_4 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_4_io_en),
    .io_configuration(Multiplexer_4_io_configuration),
    .io_inputs_3(Multiplexer_4_io_inputs_3),
    .io_inputs_2(Multiplexer_4_io_inputs_2),
    .io_inputs_1(Multiplexer_4_io_inputs_1),
    .io_inputs_0(Multiplexer_4_io_inputs_0),
    .io_outs_0(Multiplexer_4_io_outs_0)
  );
  Multiplexer Multiplexer_5 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_5_io_en),
    .io_configuration(Multiplexer_5_io_configuration),
    .io_inputs_3(Multiplexer_5_io_inputs_3),
    .io_inputs_2(Multiplexer_5_io_inputs_2),
    .io_inputs_1(Multiplexer_5_io_inputs_1),
    .io_inputs_0(Multiplexer_5_io_inputs_0),
    .io_outs_0(Multiplexer_5_io_outs_0)
  );
  Multiplexer Multiplexer_6 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_6_io_en),
    .io_configuration(Multiplexer_6_io_configuration),
    .io_inputs_3(Multiplexer_6_io_inputs_3),
    .io_inputs_2(Multiplexer_6_io_inputs_2),
    .io_inputs_1(Multiplexer_6_io_inputs_1),
    .io_inputs_0(Multiplexer_6_io_inputs_0),
    .io_outs_0(Multiplexer_6_io_outs_0)
  );
  Multiplexer Multiplexer_7 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_7_io_en),
    .io_configuration(Multiplexer_7_io_configuration),
    .io_inputs_3(Multiplexer_7_io_inputs_3),
    .io_inputs_2(Multiplexer_7_io_inputs_2),
    .io_inputs_1(Multiplexer_7_io_inputs_1),
    .io_inputs_0(Multiplexer_7_io_inputs_0),
    .io_outs_0(Multiplexer_7_io_outs_0)
  );
  Multiplexer_8 Multiplexer_8 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_8_io_en),
    .io_configuration(Multiplexer_8_io_configuration),
    .io_inputs_7(Multiplexer_8_io_inputs_7),
    .io_inputs_6(Multiplexer_8_io_inputs_6),
    .io_inputs_5(Multiplexer_8_io_inputs_5),
    .io_inputs_4(Multiplexer_8_io_inputs_4),
    .io_inputs_3(Multiplexer_8_io_inputs_3),
    .io_inputs_2(Multiplexer_8_io_inputs_2),
    .io_inputs_1(Multiplexer_8_io_inputs_1),
    .io_inputs_0(Multiplexer_8_io_inputs_0),
    .io_outs_0(Multiplexer_8_io_outs_0)
  );
  Multiplexer_9 Multiplexer_9 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_9_io_en),
    .io_configuration(Multiplexer_9_io_configuration),
    .io_inputs_6(Multiplexer_9_io_inputs_6),
    .io_inputs_5(Multiplexer_9_io_inputs_5),
    .io_inputs_4(Multiplexer_9_io_inputs_4),
    .io_inputs_3(Multiplexer_9_io_inputs_3),
    .io_inputs_2(Multiplexer_9_io_inputs_2),
    .io_inputs_1(Multiplexer_9_io_inputs_1),
    .io_inputs_0(Multiplexer_9_io_inputs_0),
    .io_outs_0(Multiplexer_9_io_outs_0)
  );
  Multiplexer_8 Multiplexer_10 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_10_io_en),
    .io_configuration(Multiplexer_10_io_configuration),
    .io_inputs_7(Multiplexer_10_io_inputs_7),
    .io_inputs_6(Multiplexer_10_io_inputs_6),
    .io_inputs_5(Multiplexer_10_io_inputs_5),
    .io_inputs_4(Multiplexer_10_io_inputs_4),
    .io_inputs_3(Multiplexer_10_io_inputs_3),
    .io_inputs_2(Multiplexer_10_io_inputs_2),
    .io_inputs_1(Multiplexer_10_io_inputs_1),
    .io_inputs_0(Multiplexer_10_io_inputs_0),
    .io_outs_0(Multiplexer_10_io_outs_0)
  );
  Multiplexer_9 Multiplexer_11 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_11_io_en),
    .io_configuration(Multiplexer_11_io_configuration),
    .io_inputs_6(Multiplexer_11_io_inputs_6),
    .io_inputs_5(Multiplexer_11_io_inputs_5),
    .io_inputs_4(Multiplexer_11_io_inputs_4),
    .io_inputs_3(Multiplexer_11_io_inputs_3),
    .io_inputs_2(Multiplexer_11_io_inputs_2),
    .io_inputs_1(Multiplexer_11_io_inputs_1),
    .io_inputs_0(Multiplexer_11_io_inputs_0),
    .io_outs_0(Multiplexer_11_io_outs_0)
  );
  Multiplexer_8 Multiplexer_12 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_12_io_en),
    .io_configuration(Multiplexer_12_io_configuration),
    .io_inputs_7(Multiplexer_12_io_inputs_7),
    .io_inputs_6(Multiplexer_12_io_inputs_6),
    .io_inputs_5(Multiplexer_12_io_inputs_5),
    .io_inputs_4(Multiplexer_12_io_inputs_4),
    .io_inputs_3(Multiplexer_12_io_inputs_3),
    .io_inputs_2(Multiplexer_12_io_inputs_2),
    .io_inputs_1(Multiplexer_12_io_inputs_1),
    .io_inputs_0(Multiplexer_12_io_inputs_0),
    .io_outs_0(Multiplexer_12_io_outs_0)
  );
  Multiplexer_9 Multiplexer_13 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_13_io_en),
    .io_configuration(Multiplexer_13_io_configuration),
    .io_inputs_6(Multiplexer_13_io_inputs_6),
    .io_inputs_5(Multiplexer_13_io_inputs_5),
    .io_inputs_4(Multiplexer_13_io_inputs_4),
    .io_inputs_3(Multiplexer_13_io_inputs_3),
    .io_inputs_2(Multiplexer_13_io_inputs_2),
    .io_inputs_1(Multiplexer_13_io_inputs_1),
    .io_inputs_0(Multiplexer_13_io_inputs_0),
    .io_outs_0(Multiplexer_13_io_outs_0)
  );
  Multiplexer_8 Multiplexer_14 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_14_io_en),
    .io_configuration(Multiplexer_14_io_configuration),
    .io_inputs_7(Multiplexer_14_io_inputs_7),
    .io_inputs_6(Multiplexer_14_io_inputs_6),
    .io_inputs_5(Multiplexer_14_io_inputs_5),
    .io_inputs_4(Multiplexer_14_io_inputs_4),
    .io_inputs_3(Multiplexer_14_io_inputs_3),
    .io_inputs_2(Multiplexer_14_io_inputs_2),
    .io_inputs_1(Multiplexer_14_io_inputs_1),
    .io_inputs_0(Multiplexer_14_io_inputs_0),
    .io_outs_0(Multiplexer_14_io_outs_0)
  );
  Multiplexer_9 Multiplexer_15 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_15_io_en),
    .io_configuration(Multiplexer_15_io_configuration),
    .io_inputs_6(Multiplexer_15_io_inputs_6),
    .io_inputs_5(Multiplexer_15_io_inputs_5),
    .io_inputs_4(Multiplexer_15_io_inputs_4),
    .io_inputs_3(Multiplexer_15_io_inputs_3),
    .io_inputs_2(Multiplexer_15_io_inputs_2),
    .io_inputs_1(Multiplexer_15_io_inputs_1),
    .io_inputs_0(Multiplexer_15_io_inputs_0),
    .io_outs_0(Multiplexer_15_io_outs_0)
  );
  Multiplexer_9 Multiplexer_16 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_16_io_en),
    .io_configuration(Multiplexer_16_io_configuration),
    .io_inputs_6(Multiplexer_16_io_inputs_6),
    .io_inputs_5(Multiplexer_16_io_inputs_5),
    .io_inputs_4(Multiplexer_16_io_inputs_4),
    .io_inputs_3(Multiplexer_16_io_inputs_3),
    .io_inputs_2(Multiplexer_16_io_inputs_2),
    .io_inputs_1(Multiplexer_16_io_inputs_1),
    .io_inputs_0(Multiplexer_16_io_inputs_0),
    .io_outs_0(Multiplexer_16_io_outs_0)
  );
  Multiplexer_17 Multiplexer_17 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_17_io_en),
    .io_configuration(Multiplexer_17_io_configuration),
    .io_inputs_5(Multiplexer_17_io_inputs_5),
    .io_inputs_4(Multiplexer_17_io_inputs_4),
    .io_inputs_3(Multiplexer_17_io_inputs_3),
    .io_inputs_2(Multiplexer_17_io_inputs_2),
    .io_inputs_1(Multiplexer_17_io_inputs_1),
    .io_inputs_0(Multiplexer_17_io_inputs_0),
    .io_outs_0(Multiplexer_17_io_outs_0)
  );
  Multiplexer_9 Multiplexer_18 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_18_io_en),
    .io_configuration(Multiplexer_18_io_configuration),
    .io_inputs_6(Multiplexer_18_io_inputs_6),
    .io_inputs_5(Multiplexer_18_io_inputs_5),
    .io_inputs_4(Multiplexer_18_io_inputs_4),
    .io_inputs_3(Multiplexer_18_io_inputs_3),
    .io_inputs_2(Multiplexer_18_io_inputs_2),
    .io_inputs_1(Multiplexer_18_io_inputs_1),
    .io_inputs_0(Multiplexer_18_io_inputs_0),
    .io_outs_0(Multiplexer_18_io_outs_0)
  );
  Multiplexer_17 Multiplexer_19 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_19_io_en),
    .io_configuration(Multiplexer_19_io_configuration),
    .io_inputs_5(Multiplexer_19_io_inputs_5),
    .io_inputs_4(Multiplexer_19_io_inputs_4),
    .io_inputs_3(Multiplexer_19_io_inputs_3),
    .io_inputs_2(Multiplexer_19_io_inputs_2),
    .io_inputs_1(Multiplexer_19_io_inputs_1),
    .io_inputs_0(Multiplexer_19_io_inputs_0),
    .io_outs_0(Multiplexer_19_io_outs_0)
  );
  Multiplexer_9 Multiplexer_20 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_20_io_en),
    .io_configuration(Multiplexer_20_io_configuration),
    .io_inputs_6(Multiplexer_20_io_inputs_6),
    .io_inputs_5(Multiplexer_20_io_inputs_5),
    .io_inputs_4(Multiplexer_20_io_inputs_4),
    .io_inputs_3(Multiplexer_20_io_inputs_3),
    .io_inputs_2(Multiplexer_20_io_inputs_2),
    .io_inputs_1(Multiplexer_20_io_inputs_1),
    .io_inputs_0(Multiplexer_20_io_inputs_0),
    .io_outs_0(Multiplexer_20_io_outs_0)
  );
  Multiplexer_17 Multiplexer_21 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_21_io_en),
    .io_configuration(Multiplexer_21_io_configuration),
    .io_inputs_5(Multiplexer_21_io_inputs_5),
    .io_inputs_4(Multiplexer_21_io_inputs_4),
    .io_inputs_3(Multiplexer_21_io_inputs_3),
    .io_inputs_2(Multiplexer_21_io_inputs_2),
    .io_inputs_1(Multiplexer_21_io_inputs_1),
    .io_inputs_0(Multiplexer_21_io_inputs_0),
    .io_outs_0(Multiplexer_21_io_outs_0)
  );
  Multiplexer_9 Multiplexer_22 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_22_io_en),
    .io_configuration(Multiplexer_22_io_configuration),
    .io_inputs_6(Multiplexer_22_io_inputs_6),
    .io_inputs_5(Multiplexer_22_io_inputs_5),
    .io_inputs_4(Multiplexer_22_io_inputs_4),
    .io_inputs_3(Multiplexer_22_io_inputs_3),
    .io_inputs_2(Multiplexer_22_io_inputs_2),
    .io_inputs_1(Multiplexer_22_io_inputs_1),
    .io_inputs_0(Multiplexer_22_io_inputs_0),
    .io_outs_0(Multiplexer_22_io_outs_0)
  );
  Multiplexer_17 Multiplexer_23 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_23_io_en),
    .io_configuration(Multiplexer_23_io_configuration),
    .io_inputs_5(Multiplexer_23_io_inputs_5),
    .io_inputs_4(Multiplexer_23_io_inputs_4),
    .io_inputs_3(Multiplexer_23_io_inputs_3),
    .io_inputs_2(Multiplexer_23_io_inputs_2),
    .io_inputs_1(Multiplexer_23_io_inputs_1),
    .io_inputs_0(Multiplexer_23_io_inputs_0),
    .io_outs_0(Multiplexer_23_io_outs_0)
  );
  Multiplexer_9 Multiplexer_24 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_24_io_en),
    .io_configuration(Multiplexer_24_io_configuration),
    .io_inputs_6(Multiplexer_24_io_inputs_6),
    .io_inputs_5(Multiplexer_24_io_inputs_5),
    .io_inputs_4(Multiplexer_24_io_inputs_4),
    .io_inputs_3(Multiplexer_24_io_inputs_3),
    .io_inputs_2(Multiplexer_24_io_inputs_2),
    .io_inputs_1(Multiplexer_24_io_inputs_1),
    .io_inputs_0(Multiplexer_24_io_inputs_0),
    .io_outs_0(Multiplexer_24_io_outs_0)
  );
  Multiplexer_17 Multiplexer_25 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_25_io_en),
    .io_configuration(Multiplexer_25_io_configuration),
    .io_inputs_5(Multiplexer_25_io_inputs_5),
    .io_inputs_4(Multiplexer_25_io_inputs_4),
    .io_inputs_3(Multiplexer_25_io_inputs_3),
    .io_inputs_2(Multiplexer_25_io_inputs_2),
    .io_inputs_1(Multiplexer_25_io_inputs_1),
    .io_inputs_0(Multiplexer_25_io_inputs_0),
    .io_outs_0(Multiplexer_25_io_outs_0)
  );
  Multiplexer_9 Multiplexer_26 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_26_io_en),
    .io_configuration(Multiplexer_26_io_configuration),
    .io_inputs_6(Multiplexer_26_io_inputs_6),
    .io_inputs_5(Multiplexer_26_io_inputs_5),
    .io_inputs_4(Multiplexer_26_io_inputs_4),
    .io_inputs_3(Multiplexer_26_io_inputs_3),
    .io_inputs_2(Multiplexer_26_io_inputs_2),
    .io_inputs_1(Multiplexer_26_io_inputs_1),
    .io_inputs_0(Multiplexer_26_io_inputs_0),
    .io_outs_0(Multiplexer_26_io_outs_0)
  );
  Multiplexer_17 Multiplexer_27 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_27_io_en),
    .io_configuration(Multiplexer_27_io_configuration),
    .io_inputs_5(Multiplexer_27_io_inputs_5),
    .io_inputs_4(Multiplexer_27_io_inputs_4),
    .io_inputs_3(Multiplexer_27_io_inputs_3),
    .io_inputs_2(Multiplexer_27_io_inputs_2),
    .io_inputs_1(Multiplexer_27_io_inputs_1),
    .io_inputs_0(Multiplexer_27_io_inputs_0),
    .io_outs_0(Multiplexer_27_io_outs_0)
  );
  Multiplexer_9 Multiplexer_28 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_28_io_en),
    .io_configuration(Multiplexer_28_io_configuration),
    .io_inputs_6(Multiplexer_28_io_inputs_6),
    .io_inputs_5(Multiplexer_28_io_inputs_5),
    .io_inputs_4(Multiplexer_28_io_inputs_4),
    .io_inputs_3(Multiplexer_28_io_inputs_3),
    .io_inputs_2(Multiplexer_28_io_inputs_2),
    .io_inputs_1(Multiplexer_28_io_inputs_1),
    .io_inputs_0(Multiplexer_28_io_inputs_0),
    .io_outs_0(Multiplexer_28_io_outs_0)
  );
  Multiplexer_17 Multiplexer_29 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_29_io_en),
    .io_configuration(Multiplexer_29_io_configuration),
    .io_inputs_5(Multiplexer_29_io_inputs_5),
    .io_inputs_4(Multiplexer_29_io_inputs_4),
    .io_inputs_3(Multiplexer_29_io_inputs_3),
    .io_inputs_2(Multiplexer_29_io_inputs_2),
    .io_inputs_1(Multiplexer_29_io_inputs_1),
    .io_inputs_0(Multiplexer_29_io_inputs_0),
    .io_outs_0(Multiplexer_29_io_outs_0)
  );
  Multiplexer_9 Multiplexer_30 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_30_io_en),
    .io_configuration(Multiplexer_30_io_configuration),
    .io_inputs_6(Multiplexer_30_io_inputs_6),
    .io_inputs_5(Multiplexer_30_io_inputs_5),
    .io_inputs_4(Multiplexer_30_io_inputs_4),
    .io_inputs_3(Multiplexer_30_io_inputs_3),
    .io_inputs_2(Multiplexer_30_io_inputs_2),
    .io_inputs_1(Multiplexer_30_io_inputs_1),
    .io_inputs_0(Multiplexer_30_io_inputs_0),
    .io_outs_0(Multiplexer_30_io_outs_0)
  );
  Multiplexer_17 Multiplexer_31 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_31_io_en),
    .io_configuration(Multiplexer_31_io_configuration),
    .io_inputs_5(Multiplexer_31_io_inputs_5),
    .io_inputs_4(Multiplexer_31_io_inputs_4),
    .io_inputs_3(Multiplexer_31_io_inputs_3),
    .io_inputs_2(Multiplexer_31_io_inputs_2),
    .io_inputs_1(Multiplexer_31_io_inputs_1),
    .io_inputs_0(Multiplexer_31_io_inputs_0),
    .io_outs_0(Multiplexer_31_io_outs_0)
  );
  Multiplexer_9 Multiplexer_32 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_32_io_en),
    .io_configuration(Multiplexer_32_io_configuration),
    .io_inputs_6(Multiplexer_32_io_inputs_6),
    .io_inputs_5(Multiplexer_32_io_inputs_5),
    .io_inputs_4(Multiplexer_32_io_inputs_4),
    .io_inputs_3(Multiplexer_32_io_inputs_3),
    .io_inputs_2(Multiplexer_32_io_inputs_2),
    .io_inputs_1(Multiplexer_32_io_inputs_1),
    .io_inputs_0(Multiplexer_32_io_inputs_0),
    .io_outs_0(Multiplexer_32_io_outs_0)
  );
  Multiplexer_17 Multiplexer_33 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_33_io_en),
    .io_configuration(Multiplexer_33_io_configuration),
    .io_inputs_5(Multiplexer_33_io_inputs_5),
    .io_inputs_4(Multiplexer_33_io_inputs_4),
    .io_inputs_3(Multiplexer_33_io_inputs_3),
    .io_inputs_2(Multiplexer_33_io_inputs_2),
    .io_inputs_1(Multiplexer_33_io_inputs_1),
    .io_inputs_0(Multiplexer_33_io_inputs_0),
    .io_outs_0(Multiplexer_33_io_outs_0)
  );
  Multiplexer_9 Multiplexer_34 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_34_io_en),
    .io_configuration(Multiplexer_34_io_configuration),
    .io_inputs_6(Multiplexer_34_io_inputs_6),
    .io_inputs_5(Multiplexer_34_io_inputs_5),
    .io_inputs_4(Multiplexer_34_io_inputs_4),
    .io_inputs_3(Multiplexer_34_io_inputs_3),
    .io_inputs_2(Multiplexer_34_io_inputs_2),
    .io_inputs_1(Multiplexer_34_io_inputs_1),
    .io_inputs_0(Multiplexer_34_io_inputs_0),
    .io_outs_0(Multiplexer_34_io_outs_0)
  );
  Multiplexer_17 Multiplexer_35 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_35_io_en),
    .io_configuration(Multiplexer_35_io_configuration),
    .io_inputs_5(Multiplexer_35_io_inputs_5),
    .io_inputs_4(Multiplexer_35_io_inputs_4),
    .io_inputs_3(Multiplexer_35_io_inputs_3),
    .io_inputs_2(Multiplexer_35_io_inputs_2),
    .io_inputs_1(Multiplexer_35_io_inputs_1),
    .io_inputs_0(Multiplexer_35_io_inputs_0),
    .io_outs_0(Multiplexer_35_io_outs_0)
  );
  Multiplexer_9 Multiplexer_36 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_36_io_en),
    .io_configuration(Multiplexer_36_io_configuration),
    .io_inputs_6(Multiplexer_36_io_inputs_6),
    .io_inputs_5(Multiplexer_36_io_inputs_5),
    .io_inputs_4(Multiplexer_36_io_inputs_4),
    .io_inputs_3(Multiplexer_36_io_inputs_3),
    .io_inputs_2(Multiplexer_36_io_inputs_2),
    .io_inputs_1(Multiplexer_36_io_inputs_1),
    .io_inputs_0(Multiplexer_36_io_inputs_0),
    .io_outs_0(Multiplexer_36_io_outs_0)
  );
  Multiplexer_17 Multiplexer_37 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_37_io_en),
    .io_configuration(Multiplexer_37_io_configuration),
    .io_inputs_5(Multiplexer_37_io_inputs_5),
    .io_inputs_4(Multiplexer_37_io_inputs_4),
    .io_inputs_3(Multiplexer_37_io_inputs_3),
    .io_inputs_2(Multiplexer_37_io_inputs_2),
    .io_inputs_1(Multiplexer_37_io_inputs_1),
    .io_inputs_0(Multiplexer_37_io_inputs_0),
    .io_outs_0(Multiplexer_37_io_outs_0)
  );
  Multiplexer_9 Multiplexer_38 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_38_io_en),
    .io_configuration(Multiplexer_38_io_configuration),
    .io_inputs_6(Multiplexer_38_io_inputs_6),
    .io_inputs_5(Multiplexer_38_io_inputs_5),
    .io_inputs_4(Multiplexer_38_io_inputs_4),
    .io_inputs_3(Multiplexer_38_io_inputs_3),
    .io_inputs_2(Multiplexer_38_io_inputs_2),
    .io_inputs_1(Multiplexer_38_io_inputs_1),
    .io_inputs_0(Multiplexer_38_io_inputs_0),
    .io_outs_0(Multiplexer_38_io_outs_0)
  );
  Multiplexer_17 Multiplexer_39 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_39_io_en),
    .io_configuration(Multiplexer_39_io_configuration),
    .io_inputs_5(Multiplexer_39_io_inputs_5),
    .io_inputs_4(Multiplexer_39_io_inputs_4),
    .io_inputs_3(Multiplexer_39_io_inputs_3),
    .io_inputs_2(Multiplexer_39_io_inputs_2),
    .io_inputs_1(Multiplexer_39_io_inputs_1),
    .io_inputs_0(Multiplexer_39_io_inputs_0),
    .io_outs_0(Multiplexer_39_io_outs_0)
  );
  Multiplexer Multiplexer_40 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_40_io_en),
    .io_configuration(Multiplexer_40_io_configuration),
    .io_inputs_3(Multiplexer_40_io_inputs_3),
    .io_inputs_2(Multiplexer_40_io_inputs_2),
    .io_inputs_1(Multiplexer_40_io_inputs_1),
    .io_inputs_0(Multiplexer_40_io_inputs_0),
    .io_outs_0(Multiplexer_40_io_outs_0)
  );
  Multiplexer Multiplexer_41 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_41_io_en),
    .io_configuration(Multiplexer_41_io_configuration),
    .io_inputs_3(Multiplexer_41_io_inputs_3),
    .io_inputs_2(Multiplexer_41_io_inputs_2),
    .io_inputs_1(Multiplexer_41_io_inputs_1),
    .io_inputs_0(Multiplexer_41_io_inputs_0),
    .io_outs_0(Multiplexer_41_io_outs_0)
  );
  Multiplexer Multiplexer_42 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_42_io_en),
    .io_configuration(Multiplexer_42_io_configuration),
    .io_inputs_3(Multiplexer_42_io_inputs_3),
    .io_inputs_2(Multiplexer_42_io_inputs_2),
    .io_inputs_1(Multiplexer_42_io_inputs_1),
    .io_inputs_0(Multiplexer_42_io_inputs_0),
    .io_outs_0(Multiplexer_42_io_outs_0)
  );
  Multiplexer Multiplexer_43 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_43_io_en),
    .io_configuration(Multiplexer_43_io_configuration),
    .io_inputs_3(Multiplexer_43_io_inputs_3),
    .io_inputs_2(Multiplexer_43_io_inputs_2),
    .io_inputs_1(Multiplexer_43_io_inputs_1),
    .io_inputs_0(Multiplexer_43_io_inputs_0),
    .io_outs_0(Multiplexer_43_io_outs_0)
  );
  Multiplexer Multiplexer_44 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_44_io_en),
    .io_configuration(Multiplexer_44_io_configuration),
    .io_inputs_3(Multiplexer_44_io_inputs_3),
    .io_inputs_2(Multiplexer_44_io_inputs_2),
    .io_inputs_1(Multiplexer_44_io_inputs_1),
    .io_inputs_0(Multiplexer_44_io_inputs_0),
    .io_outs_0(Multiplexer_44_io_outs_0)
  );
  Multiplexer Multiplexer_45 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_45_io_en),
    .io_configuration(Multiplexer_45_io_configuration),
    .io_inputs_3(Multiplexer_45_io_inputs_3),
    .io_inputs_2(Multiplexer_45_io_inputs_2),
    .io_inputs_1(Multiplexer_45_io_inputs_1),
    .io_inputs_0(Multiplexer_45_io_inputs_0),
    .io_outs_0(Multiplexer_45_io_outs_0)
  );
  Multiplexer Multiplexer_46 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_46_io_en),
    .io_configuration(Multiplexer_46_io_configuration),
    .io_inputs_3(Multiplexer_46_io_inputs_3),
    .io_inputs_2(Multiplexer_46_io_inputs_2),
    .io_inputs_1(Multiplexer_46_io_inputs_1),
    .io_inputs_0(Multiplexer_46_io_inputs_0),
    .io_outs_0(Multiplexer_46_io_outs_0)
  );
  Multiplexer Multiplexer_47 ( // @[TopModule.scala 154:11]
    .io_en(Multiplexer_47_io_en),
    .io_configuration(Multiplexer_47_io_configuration),
    .io_inputs_3(Multiplexer_47_io_inputs_3),
    .io_inputs_2(Multiplexer_47_io_inputs_2),
    .io_inputs_1(Multiplexer_47_io_inputs_1),
    .io_inputs_0(Multiplexer_47_io_inputs_0),
    .io_outs_0(Multiplexer_47_io_outs_0)
  );
  ConstUnit ConstUnit ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_io_en),
    .io_configuration(ConstUnit_io_configuration),
    .io_outs_0(ConstUnit_io_outs_0)
  );
  ConstUnit ConstUnit_1 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_1_io_en),
    .io_configuration(ConstUnit_1_io_configuration),
    .io_outs_0(ConstUnit_1_io_outs_0)
  );
  ConstUnit ConstUnit_2 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_2_io_en),
    .io_configuration(ConstUnit_2_io_configuration),
    .io_outs_0(ConstUnit_2_io_outs_0)
  );
  ConstUnit ConstUnit_3 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_3_io_en),
    .io_configuration(ConstUnit_3_io_configuration),
    .io_outs_0(ConstUnit_3_io_outs_0)
  );
  ConstUnit ConstUnit_4 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_4_io_en),
    .io_configuration(ConstUnit_4_io_configuration),
    .io_outs_0(ConstUnit_4_io_outs_0)
  );
  ConstUnit ConstUnit_5 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_5_io_en),
    .io_configuration(ConstUnit_5_io_configuration),
    .io_outs_0(ConstUnit_5_io_outs_0)
  );
  ConstUnit ConstUnit_6 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_6_io_en),
    .io_configuration(ConstUnit_6_io_configuration),
    .io_outs_0(ConstUnit_6_io_outs_0)
  );
  ConstUnit ConstUnit_7 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_7_io_en),
    .io_configuration(ConstUnit_7_io_configuration),
    .io_outs_0(ConstUnit_7_io_outs_0)
  );
  ConstUnit ConstUnit_8 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_8_io_en),
    .io_configuration(ConstUnit_8_io_configuration),
    .io_outs_0(ConstUnit_8_io_outs_0)
  );
  ConstUnit ConstUnit_9 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_9_io_en),
    .io_configuration(ConstUnit_9_io_configuration),
    .io_outs_0(ConstUnit_9_io_outs_0)
  );
  ConstUnit ConstUnit_10 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_10_io_en),
    .io_configuration(ConstUnit_10_io_configuration),
    .io_outs_0(ConstUnit_10_io_outs_0)
  );
  ConstUnit ConstUnit_11 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_11_io_en),
    .io_configuration(ConstUnit_11_io_configuration),
    .io_outs_0(ConstUnit_11_io_outs_0)
  );
  ConstUnit ConstUnit_12 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_12_io_en),
    .io_configuration(ConstUnit_12_io_configuration),
    .io_outs_0(ConstUnit_12_io_outs_0)
  );
  ConstUnit ConstUnit_13 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_13_io_en),
    .io_configuration(ConstUnit_13_io_configuration),
    .io_outs_0(ConstUnit_13_io_outs_0)
  );
  ConstUnit ConstUnit_14 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_14_io_en),
    .io_configuration(ConstUnit_14_io_configuration),
    .io_outs_0(ConstUnit_14_io_outs_0)
  );
  ConstUnit ConstUnit_15 ( // @[TopModule.scala 163:21]
    .io_en(ConstUnit_15_io_en),
    .io_configuration(ConstUnit_15_io_configuration),
    .io_outs_0(ConstUnit_15_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit ( // @[TopModule.scala 171:21]
    .clock(LoadStoreUnit_clock),
    .reset(LoadStoreUnit_reset),
    .io_configuration(LoadStoreUnit_io_configuration),
    .io_en(LoadStoreUnit_io_en),
    .io_skewing(LoadStoreUnit_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_io_streamIn_bits),
    .io_len(LoadStoreUnit_io_len),
    .io_streamOut_ready(LoadStoreUnit_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_io_streamOut_bits),
    .io_base(LoadStoreUnit_io_base),
    .io_start(LoadStoreUnit_io_start),
    .io_enqEn(LoadStoreUnit_io_enqEn),
    .io_deqEn(LoadStoreUnit_io_deqEn),
    .io_idle(LoadStoreUnit_io_idle),
    .io_inputs_1(LoadStoreUnit_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_io_inputs_0),
    .io_outs_0(LoadStoreUnit_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_1 ( // @[TopModule.scala 171:21]
    .clock(LoadStoreUnit_1_clock),
    .reset(LoadStoreUnit_1_reset),
    .io_configuration(LoadStoreUnit_1_io_configuration),
    .io_en(LoadStoreUnit_1_io_en),
    .io_skewing(LoadStoreUnit_1_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_1_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_1_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_1_io_streamIn_bits),
    .io_len(LoadStoreUnit_1_io_len),
    .io_streamOut_ready(LoadStoreUnit_1_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_1_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_1_io_streamOut_bits),
    .io_base(LoadStoreUnit_1_io_base),
    .io_start(LoadStoreUnit_1_io_start),
    .io_enqEn(LoadStoreUnit_1_io_enqEn),
    .io_deqEn(LoadStoreUnit_1_io_deqEn),
    .io_idle(LoadStoreUnit_1_io_idle),
    .io_inputs_1(LoadStoreUnit_1_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_1_io_inputs_0),
    .io_outs_0(LoadStoreUnit_1_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_2 ( // @[TopModule.scala 171:21]
    .clock(LoadStoreUnit_2_clock),
    .reset(LoadStoreUnit_2_reset),
    .io_configuration(LoadStoreUnit_2_io_configuration),
    .io_en(LoadStoreUnit_2_io_en),
    .io_skewing(LoadStoreUnit_2_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_2_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_2_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_2_io_streamIn_bits),
    .io_len(LoadStoreUnit_2_io_len),
    .io_streamOut_ready(LoadStoreUnit_2_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_2_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_2_io_streamOut_bits),
    .io_base(LoadStoreUnit_2_io_base),
    .io_start(LoadStoreUnit_2_io_start),
    .io_enqEn(LoadStoreUnit_2_io_enqEn),
    .io_deqEn(LoadStoreUnit_2_io_deqEn),
    .io_idle(LoadStoreUnit_2_io_idle),
    .io_inputs_1(LoadStoreUnit_2_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_2_io_inputs_0),
    .io_outs_0(LoadStoreUnit_2_io_outs_0)
  );
  LoadStoreUnit LoadStoreUnit_3 ( // @[TopModule.scala 171:21]
    .clock(LoadStoreUnit_3_clock),
    .reset(LoadStoreUnit_3_reset),
    .io_configuration(LoadStoreUnit_3_io_configuration),
    .io_en(LoadStoreUnit_3_io_en),
    .io_skewing(LoadStoreUnit_3_io_skewing),
    .io_streamIn_ready(LoadStoreUnit_3_io_streamIn_ready),
    .io_streamIn_valid(LoadStoreUnit_3_io_streamIn_valid),
    .io_streamIn_bits(LoadStoreUnit_3_io_streamIn_bits),
    .io_len(LoadStoreUnit_3_io_len),
    .io_streamOut_ready(LoadStoreUnit_3_io_streamOut_ready),
    .io_streamOut_valid(LoadStoreUnit_3_io_streamOut_valid),
    .io_streamOut_bits(LoadStoreUnit_3_io_streamOut_bits),
    .io_base(LoadStoreUnit_3_io_base),
    .io_start(LoadStoreUnit_3_io_start),
    .io_enqEn(LoadStoreUnit_3_io_enqEn),
    .io_deqEn(LoadStoreUnit_3_io_deqEn),
    .io_idle(LoadStoreUnit_3_io_idle),
    .io_inputs_1(LoadStoreUnit_3_io_inputs_1),
    .io_inputs_0(LoadStoreUnit_3_io_inputs_0),
    .io_outs_0(LoadStoreUnit_3_io_outs_0)
  );
  MultiIIScheduleController MultiIIScheduleController_16 ( // @[TopModule.scala 172:78]
    .clock(MultiIIScheduleController_16_clock),
    .reset(MultiIIScheduleController_16_reset),
    .io_en(MultiIIScheduleController_16_io_en),
    .io_schedules_0(MultiIIScheduleController_16_io_schedules_0),
    .io_II(MultiIIScheduleController_16_io_II),
    .io_valid(MultiIIScheduleController_16_io_valid),
    .io_skewing(MultiIIScheduleController_16_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_17 ( // @[TopModule.scala 172:78]
    .clock(MultiIIScheduleController_17_clock),
    .reset(MultiIIScheduleController_17_reset),
    .io_en(MultiIIScheduleController_17_io_en),
    .io_schedules_0(MultiIIScheduleController_17_io_schedules_0),
    .io_II(MultiIIScheduleController_17_io_II),
    .io_valid(MultiIIScheduleController_17_io_valid),
    .io_skewing(MultiIIScheduleController_17_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_18 ( // @[TopModule.scala 172:78]
    .clock(MultiIIScheduleController_18_clock),
    .reset(MultiIIScheduleController_18_reset),
    .io_en(MultiIIScheduleController_18_io_en),
    .io_schedules_0(MultiIIScheduleController_18_io_schedules_0),
    .io_II(MultiIIScheduleController_18_io_II),
    .io_valid(MultiIIScheduleController_18_io_valid),
    .io_skewing(MultiIIScheduleController_18_io_skewing)
  );
  MultiIIScheduleController MultiIIScheduleController_19 ( // @[TopModule.scala 172:78]
    .clock(MultiIIScheduleController_19_clock),
    .reset(MultiIIScheduleController_19_reset),
    .io_en(MultiIIScheduleController_19_io_en),
    .io_schedules_0(MultiIIScheduleController_19_io_schedules_0),
    .io_II(MultiIIScheduleController_19_io_II),
    .io_valid(MultiIIScheduleController_19_io_valid),
    .io_skewing(MultiIIScheduleController_19_io_skewing)
  );
  ConfigController configController ( // @[TopModule.scala 219:32]
    .clock(configController_clock),
    .reset(configController_reset),
    .io_en(configController_io_en),
    .io_II(configController_io_II),
    .io_outConfig(configController_io_outConfig)
  );
  Dispatch_14 dispatchs_0 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_0_io_en),
    .io_configuration(dispatchs_0_io_configuration),
    .io_outs_3(dispatchs_0_io_outs_3),
    .io_outs_2(dispatchs_0_io_outs_2),
    .io_outs_1(dispatchs_0_io_outs_1),
    .io_outs_0(dispatchs_0_io_outs_0)
  );
  Dispatch_15 dispatchs_1 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_1_io_en),
    .io_configuration(dispatchs_1_io_configuration),
    .io_outs_4(dispatchs_1_io_outs_4),
    .io_outs_3(dispatchs_1_io_outs_3),
    .io_outs_2(dispatchs_1_io_outs_2),
    .io_outs_1(dispatchs_1_io_outs_1),
    .io_outs_0(dispatchs_1_io_outs_0)
  );
  Dispatch_14 dispatchs_2 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_2_io_en),
    .io_configuration(dispatchs_2_io_configuration),
    .io_outs_3(dispatchs_2_io_outs_3),
    .io_outs_2(dispatchs_2_io_outs_2),
    .io_outs_1(dispatchs_2_io_outs_1),
    .io_outs_0(dispatchs_2_io_outs_0)
  );
  Dispatch_15 dispatchs_3 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_3_io_en),
    .io_configuration(dispatchs_3_io_configuration),
    .io_outs_4(dispatchs_3_io_outs_4),
    .io_outs_3(dispatchs_3_io_outs_3),
    .io_outs_2(dispatchs_3_io_outs_2),
    .io_outs_1(dispatchs_3_io_outs_1),
    .io_outs_0(dispatchs_3_io_outs_0)
  );
  Dispatch_15 dispatchs_4 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_4_io_en),
    .io_configuration(dispatchs_4_io_configuration),
    .io_outs_4(dispatchs_4_io_outs_4),
    .io_outs_3(dispatchs_4_io_outs_3),
    .io_outs_2(dispatchs_4_io_outs_2),
    .io_outs_1(dispatchs_4_io_outs_1),
    .io_outs_0(dispatchs_4_io_outs_0)
  );
  Dispatch_19 dispatchs_5 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_5_io_en),
    .io_configuration(dispatchs_5_io_configuration),
    .io_outs_7(dispatchs_5_io_outs_7),
    .io_outs_6(dispatchs_5_io_outs_6),
    .io_outs_5(dispatchs_5_io_outs_5),
    .io_outs_4(dispatchs_5_io_outs_4),
    .io_outs_3(dispatchs_5_io_outs_3),
    .io_outs_2(dispatchs_5_io_outs_2),
    .io_outs_1(dispatchs_5_io_outs_1),
    .io_outs_0(dispatchs_5_io_outs_0)
  );
  Dispatch_15 dispatchs_6 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_6_io_en),
    .io_configuration(dispatchs_6_io_configuration),
    .io_outs_4(dispatchs_6_io_outs_4),
    .io_outs_3(dispatchs_6_io_outs_3),
    .io_outs_2(dispatchs_6_io_outs_2),
    .io_outs_1(dispatchs_6_io_outs_1),
    .io_outs_0(dispatchs_6_io_outs_0)
  );
  Dispatch_21 dispatchs_7 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_7_io_en),
    .io_configuration(dispatchs_7_io_configuration),
    .io_outs_2(dispatchs_7_io_outs_2),
    .io_outs_1(dispatchs_7_io_outs_1),
    .io_outs_0(dispatchs_7_io_outs_0)
  );
  Dispatch_15 dispatchs_8 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_8_io_en),
    .io_configuration(dispatchs_8_io_configuration),
    .io_outs_4(dispatchs_8_io_outs_4),
    .io_outs_3(dispatchs_8_io_outs_3),
    .io_outs_2(dispatchs_8_io_outs_2),
    .io_outs_1(dispatchs_8_io_outs_1),
    .io_outs_0(dispatchs_8_io_outs_0)
  );
  Dispatch_15 dispatchs_9 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_9_io_en),
    .io_configuration(dispatchs_9_io_configuration),
    .io_outs_4(dispatchs_9_io_outs_4),
    .io_outs_3(dispatchs_9_io_outs_3),
    .io_outs_2(dispatchs_9_io_outs_2),
    .io_outs_1(dispatchs_9_io_outs_1),
    .io_outs_0(dispatchs_9_io_outs_0)
  );
  Dispatch_15 dispatchs_10 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_10_io_en),
    .io_configuration(dispatchs_10_io_configuration),
    .io_outs_4(dispatchs_10_io_outs_4),
    .io_outs_3(dispatchs_10_io_outs_3),
    .io_outs_2(dispatchs_10_io_outs_2),
    .io_outs_1(dispatchs_10_io_outs_1),
    .io_outs_0(dispatchs_10_io_outs_0)
  );
  Dispatch_21 dispatchs_11 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_11_io_en),
    .io_configuration(dispatchs_11_io_configuration),
    .io_outs_2(dispatchs_11_io_outs_2),
    .io_outs_1(dispatchs_11_io_outs_1),
    .io_outs_0(dispatchs_11_io_outs_0)
  );
  Dispatch_15 dispatchs_12 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_12_io_en),
    .io_configuration(dispatchs_12_io_configuration),
    .io_outs_4(dispatchs_12_io_outs_4),
    .io_outs_3(dispatchs_12_io_outs_3),
    .io_outs_2(dispatchs_12_io_outs_2),
    .io_outs_1(dispatchs_12_io_outs_1),
    .io_outs_0(dispatchs_12_io_outs_0)
  );
  Dispatch_14 dispatchs_13 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_13_io_en),
    .io_configuration(dispatchs_13_io_configuration),
    .io_outs_3(dispatchs_13_io_outs_3),
    .io_outs_2(dispatchs_13_io_outs_2),
    .io_outs_1(dispatchs_13_io_outs_1),
    .io_outs_0(dispatchs_13_io_outs_0)
  );
  Dispatch_21 dispatchs_14 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_14_io_en),
    .io_configuration(dispatchs_14_io_configuration),
    .io_outs_2(dispatchs_14_io_outs_2),
    .io_outs_1(dispatchs_14_io_outs_1),
    .io_outs_0(dispatchs_14_io_outs_0)
  );
  Dispatch_15 dispatchs_15 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_15_io_en),
    .io_configuration(dispatchs_15_io_configuration),
    .io_outs_4(dispatchs_15_io_outs_4),
    .io_outs_3(dispatchs_15_io_outs_3),
    .io_outs_2(dispatchs_15_io_outs_2),
    .io_outs_1(dispatchs_15_io_outs_1),
    .io_outs_0(dispatchs_15_io_outs_0)
  );
  Dispatch_30 dispatchs_16 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_16_io_en),
    .io_configuration(dispatchs_16_io_configuration),
    .io_outs_0(dispatchs_16_io_outs_0)
  );
  Dispatch_21 dispatchs_17 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_17_io_en),
    .io_configuration(dispatchs_17_io_configuration),
    .io_outs_2(dispatchs_17_io_outs_2),
    .io_outs_1(dispatchs_17_io_outs_1),
    .io_outs_0(dispatchs_17_io_outs_0)
  );
  Dispatch_15 dispatchs_18 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_18_io_en),
    .io_configuration(dispatchs_18_io_configuration),
    .io_outs_4(dispatchs_18_io_outs_4),
    .io_outs_3(dispatchs_18_io_outs_3),
    .io_outs_2(dispatchs_18_io_outs_2),
    .io_outs_1(dispatchs_18_io_outs_1),
    .io_outs_0(dispatchs_18_io_outs_0)
  );
  Dispatch_15 dispatchs_19 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_19_io_en),
    .io_configuration(dispatchs_19_io_configuration),
    .io_outs_4(dispatchs_19_io_outs_4),
    .io_outs_3(dispatchs_19_io_outs_3),
    .io_outs_2(dispatchs_19_io_outs_2),
    .io_outs_1(dispatchs_19_io_outs_1),
    .io_outs_0(dispatchs_19_io_outs_0)
  );
  Dispatch_15 dispatchs_20 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_20_io_en),
    .io_configuration(dispatchs_20_io_configuration),
    .io_outs_4(dispatchs_20_io_outs_4),
    .io_outs_3(dispatchs_20_io_outs_3),
    .io_outs_2(dispatchs_20_io_outs_2),
    .io_outs_1(dispatchs_20_io_outs_1),
    .io_outs_0(dispatchs_20_io_outs_0)
  );
  Dispatch_14 dispatchs_21 ( // @[TopModule.scala 246:26]
    .io_en(dispatchs_21_io_en),
    .io_configuration(dispatchs_21_io_configuration),
    .io_outs_3(dispatchs_21_io_outs_3),
    .io_outs_2(dispatchs_21_io_outs_2),
    .io_outs_1(dispatchs_21_io_outs_1),
    .io_outs_0(dispatchs_21_io_outs_0)
  );
  Dispatch_36 topDispatch ( // @[TopModule.scala 255:27]
    .io_en(topDispatch_io_en),
    .io_configuration(topDispatch_io_configuration),
    .io_outs_21(topDispatch_io_outs_21),
    .io_outs_20(topDispatch_io_outs_20),
    .io_outs_19(topDispatch_io_outs_19),
    .io_outs_18(topDispatch_io_outs_18),
    .io_outs_17(topDispatch_io_outs_17),
    .io_outs_16(topDispatch_io_outs_16),
    .io_outs_15(topDispatch_io_outs_15),
    .io_outs_14(topDispatch_io_outs_14),
    .io_outs_13(topDispatch_io_outs_13),
    .io_outs_12(topDispatch_io_outs_12),
    .io_outs_11(topDispatch_io_outs_11),
    .io_outs_10(topDispatch_io_outs_10),
    .io_outs_9(topDispatch_io_outs_9),
    .io_outs_8(topDispatch_io_outs_8),
    .io_outs_7(topDispatch_io_outs_7),
    .io_outs_6(topDispatch_io_outs_6),
    .io_outs_5(topDispatch_io_outs_5),
    .io_outs_4(topDispatch_io_outs_4),
    .io_outs_3(topDispatch_io_outs_3),
    .io_outs_2(topDispatch_io_outs_2),
    .io_outs_1(topDispatch_io_outs_1),
    .io_outs_0(topDispatch_io_outs_0)
  );
  assign io_streamInLSU_3_ready = LoadStoreUnit_3_io_streamIn_ready; // @[TopModule.scala 184:21]
  assign io_streamInLSU_2_ready = LoadStoreUnit_2_io_streamIn_ready; // @[TopModule.scala 184:21]
  assign io_streamInLSU_1_ready = LoadStoreUnit_1_io_streamIn_ready; // @[TopModule.scala 184:21]
  assign io_streamInLSU_0_ready = LoadStoreUnit_io_streamIn_ready; // @[TopModule.scala 184:21]
  assign io_streamOutLSU_3_valid = LoadStoreUnit_3_io_streamOut_valid; // @[TopModule.scala 185:22]
  assign io_streamOutLSU_3_bits = LoadStoreUnit_3_io_streamOut_bits; // @[TopModule.scala 185:22]
  assign io_streamOutLSU_2_valid = LoadStoreUnit_2_io_streamOut_valid; // @[TopModule.scala 185:22]
  assign io_streamOutLSU_2_bits = LoadStoreUnit_2_io_streamOut_bits; // @[TopModule.scala 185:22]
  assign io_streamOutLSU_1_valid = LoadStoreUnit_1_io_streamOut_valid; // @[TopModule.scala 185:22]
  assign io_streamOutLSU_1_bits = LoadStoreUnit_1_io_streamOut_bits; // @[TopModule.scala 185:22]
  assign io_streamOutLSU_0_valid = LoadStoreUnit_io_streamOut_valid; // @[TopModule.scala 185:22]
  assign io_streamOutLSU_0_bits = LoadStoreUnit_io_streamOut_bits; // @[TopModule.scala 185:22]
  assign io_idleLSU_0 = LoadStoreUnit_io_idle; // @[TopModule.scala 181:17]
  assign io_idleLSU_1 = LoadStoreUnit_1_io_idle; // @[TopModule.scala 181:17]
  assign io_idleLSU_2 = LoadStoreUnit_2_io_idle; // @[TopModule.scala 181:17]
  assign io_idleLSU_3 = LoadStoreUnit_3_io_idle; // @[TopModule.scala 181:17]
  assign io_outs_3 = Multiplexer_3_io_outs_0; // @[TopModule.scala 294:25]
  assign io_outs_2 = Multiplexer_2_io_outs_0; // @[TopModule.scala 294:25]
  assign io_outs_1 = Multiplexer_1_io_outs_0; // @[TopModule.scala 294:25]
  assign io_outs_0 = Multiplexer_io_outs_0; // @[TopModule.scala 294:25]
  assign scheduleDispatch_io_en = io_en; // @[TopModule.scala 121:26]
  assign Alu_clock = clock;
  assign Alu_reset = reset;
  assign Alu_io_en = MultiIIScheduleController_io_valid; // @[TopModule.scala 134:15]
  assign Alu_io_skewing = MultiIIScheduleController_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_io_configuration = dispatchs_2_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_io_inputs_1 = Multiplexer_9_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_io_inputs_0 = Multiplexer_8_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_1_clock = clock;
  assign Alu_1_reset = reset;
  assign Alu_1_io_en = MultiIIScheduleController_1_io_valid; // @[TopModule.scala 134:15]
  assign Alu_1_io_skewing = MultiIIScheduleController_1_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_1_io_configuration = dispatchs_0_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_1_io_inputs_1 = Multiplexer_11_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_1_io_inputs_0 = Multiplexer_10_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_2_clock = clock;
  assign Alu_2_reset = reset;
  assign Alu_2_io_en = MultiIIScheduleController_2_io_valid; // @[TopModule.scala 134:15]
  assign Alu_2_io_skewing = MultiIIScheduleController_2_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_2_io_configuration = dispatchs_13_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_2_io_inputs_1 = Multiplexer_13_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_2_io_inputs_0 = Multiplexer_12_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_3_clock = clock;
  assign Alu_3_reset = reset;
  assign Alu_3_io_en = MultiIIScheduleController_3_io_valid; // @[TopModule.scala 134:15]
  assign Alu_3_io_skewing = MultiIIScheduleController_3_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_3_io_configuration = dispatchs_21_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_3_io_inputs_1 = Multiplexer_15_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_3_io_inputs_0 = Multiplexer_14_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_4_clock = clock;
  assign Alu_4_reset = reset;
  assign Alu_4_io_en = MultiIIScheduleController_4_io_valid; // @[TopModule.scala 134:15]
  assign Alu_4_io_skewing = MultiIIScheduleController_4_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_4_io_configuration = dispatchs_12_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_4_io_inputs_1 = Multiplexer_17_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_4_io_inputs_0 = Multiplexer_16_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_5_clock = clock;
  assign Alu_5_reset = reset;
  assign Alu_5_io_en = MultiIIScheduleController_5_io_valid; // @[TopModule.scala 134:15]
  assign Alu_5_io_skewing = MultiIIScheduleController_5_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_5_io_configuration = dispatchs_19_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_5_io_inputs_1 = Multiplexer_19_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_5_io_inputs_0 = Multiplexer_18_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_6_clock = clock;
  assign Alu_6_reset = reset;
  assign Alu_6_io_en = MultiIIScheduleController_6_io_valid; // @[TopModule.scala 134:15]
  assign Alu_6_io_skewing = MultiIIScheduleController_6_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_6_io_configuration = dispatchs_3_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_6_io_inputs_1 = Multiplexer_21_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_6_io_inputs_0 = Multiplexer_20_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_7_clock = clock;
  assign Alu_7_reset = reset;
  assign Alu_7_io_en = MultiIIScheduleController_7_io_valid; // @[TopModule.scala 134:15]
  assign Alu_7_io_skewing = MultiIIScheduleController_7_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_7_io_configuration = dispatchs_9_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_7_io_inputs_1 = Multiplexer_23_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_7_io_inputs_0 = Multiplexer_22_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_8_clock = clock;
  assign Alu_8_reset = reset;
  assign Alu_8_io_en = MultiIIScheduleController_8_io_valid; // @[TopModule.scala 134:15]
  assign Alu_8_io_skewing = MultiIIScheduleController_8_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_8_io_configuration = dispatchs_6_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_8_io_inputs_1 = Multiplexer_25_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_8_io_inputs_0 = Multiplexer_24_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_9_clock = clock;
  assign Alu_9_reset = reset;
  assign Alu_9_io_en = MultiIIScheduleController_9_io_valid; // @[TopModule.scala 134:15]
  assign Alu_9_io_skewing = MultiIIScheduleController_9_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_9_io_configuration = dispatchs_15_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_9_io_inputs_1 = Multiplexer_27_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_9_io_inputs_0 = Multiplexer_26_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_10_clock = clock;
  assign Alu_10_reset = reset;
  assign Alu_10_io_en = MultiIIScheduleController_10_io_valid; // @[TopModule.scala 134:15]
  assign Alu_10_io_skewing = MultiIIScheduleController_10_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_10_io_configuration = dispatchs_18_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_10_io_inputs_1 = Multiplexer_29_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_10_io_inputs_0 = Multiplexer_28_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_11_clock = clock;
  assign Alu_11_reset = reset;
  assign Alu_11_io_en = MultiIIScheduleController_11_io_valid; // @[TopModule.scala 134:15]
  assign Alu_11_io_skewing = MultiIIScheduleController_11_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_11_io_configuration = dispatchs_4_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_11_io_inputs_1 = Multiplexer_31_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_11_io_inputs_0 = Multiplexer_30_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_12_clock = clock;
  assign Alu_12_reset = reset;
  assign Alu_12_io_en = MultiIIScheduleController_12_io_valid; // @[TopModule.scala 134:15]
  assign Alu_12_io_skewing = MultiIIScheduleController_12_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_12_io_configuration = dispatchs_10_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_12_io_inputs_1 = Multiplexer_33_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_12_io_inputs_0 = Multiplexer_32_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_13_clock = clock;
  assign Alu_13_reset = reset;
  assign Alu_13_io_en = MultiIIScheduleController_13_io_valid; // @[TopModule.scala 134:15]
  assign Alu_13_io_skewing = MultiIIScheduleController_13_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_13_io_configuration = dispatchs_1_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_13_io_inputs_1 = Multiplexer_35_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_13_io_inputs_0 = Multiplexer_34_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_14_clock = clock;
  assign Alu_14_reset = reset;
  assign Alu_14_io_en = MultiIIScheduleController_14_io_valid; // @[TopModule.scala 134:15]
  assign Alu_14_io_skewing = MultiIIScheduleController_14_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_14_io_configuration = dispatchs_20_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_14_io_inputs_1 = Multiplexer_37_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_14_io_inputs_0 = Multiplexer_36_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_15_clock = clock;
  assign Alu_15_reset = reset;
  assign Alu_15_io_en = MultiIIScheduleController_15_io_valid; // @[TopModule.scala 134:15]
  assign Alu_15_io_skewing = MultiIIScheduleController_15_io_skewing; // @[TopModule.scala 135:20]
  assign Alu_15_io_configuration = dispatchs_8_io_outs_0; // @[TopModule.scala 249:22]
  assign Alu_15_io_inputs_1 = Multiplexer_39_io_outs_0; // @[TopModule.scala 298:60]
  assign Alu_15_io_inputs_0 = Multiplexer_38_io_outs_0; // @[TopModule.scala 298:60]
  assign MultiIIScheduleController_clock = clock;
  assign MultiIIScheduleController_reset = reset;
  assign MultiIIScheduleController_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_1_clock = clock;
  assign MultiIIScheduleController_1_reset = reset;
  assign MultiIIScheduleController_1_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_1_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_1_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_2_clock = clock;
  assign MultiIIScheduleController_2_reset = reset;
  assign MultiIIScheduleController_2_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_2_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_2_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_3_clock = clock;
  assign MultiIIScheduleController_3_reset = reset;
  assign MultiIIScheduleController_3_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_3_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_3_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_4_clock = clock;
  assign MultiIIScheduleController_4_reset = reset;
  assign MultiIIScheduleController_4_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_4_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_4_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_5_clock = clock;
  assign MultiIIScheduleController_5_reset = reset;
  assign MultiIIScheduleController_5_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_5_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_5_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_6_clock = clock;
  assign MultiIIScheduleController_6_reset = reset;
  assign MultiIIScheduleController_6_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_6_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_6_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_7_clock = clock;
  assign MultiIIScheduleController_7_reset = reset;
  assign MultiIIScheduleController_7_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_7_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_7_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_8_clock = clock;
  assign MultiIIScheduleController_8_reset = reset;
  assign MultiIIScheduleController_8_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_8_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_8_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_9_clock = clock;
  assign MultiIIScheduleController_9_reset = reset;
  assign MultiIIScheduleController_9_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_9_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_9_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_10_clock = clock;
  assign MultiIIScheduleController_10_reset = reset;
  assign MultiIIScheduleController_10_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_10_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_10_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_11_clock = clock;
  assign MultiIIScheduleController_11_reset = reset;
  assign MultiIIScheduleController_11_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_11_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_11_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_12_clock = clock;
  assign MultiIIScheduleController_12_reset = reset;
  assign MultiIIScheduleController_12_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_12_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_12_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_13_clock = clock;
  assign MultiIIScheduleController_13_reset = reset;
  assign MultiIIScheduleController_13_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_13_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_13_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_14_clock = clock;
  assign MultiIIScheduleController_14_reset = reset;
  assign MultiIIScheduleController_14_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_14_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_14_io_II = io_II; // @[TopModule.scala 130:33]
  assign MultiIIScheduleController_15_clock = clock;
  assign MultiIIScheduleController_15_reset = reset;
  assign MultiIIScheduleController_15_io_en = io_en; // @[TopModule.scala 129:33]
  assign MultiIIScheduleController_15_io_schedules_0 = 9'h0; // @[TopModule.scala 132:45]
  assign MultiIIScheduleController_15_io_II = io_II; // @[TopModule.scala 130:33]
  assign RegisterFiles_clock = clock;
  assign RegisterFiles_reset = reset;
  assign RegisterFiles_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_io_configuration = dispatchs_16_io_outs_0; // @[TopModule.scala 249:22]
  assign RegisterFiles_io_inputs_3 = Alu_3_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_io_inputs_2 = Alu_2_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_io_inputs_1 = Alu_1_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_io_inputs_0 = Alu_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_1_clock = clock;
  assign RegisterFiles_1_reset = reset;
  assign RegisterFiles_1_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_1_io_configuration = dispatchs_12_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_1_io_inputs_0 = Alu_4_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_2_clock = clock;
  assign RegisterFiles_2_reset = reset;
  assign RegisterFiles_2_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_2_io_configuration = dispatchs_19_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_2_io_inputs_0 = Alu_5_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_3_clock = clock;
  assign RegisterFiles_3_reset = reset;
  assign RegisterFiles_3_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_3_io_configuration = dispatchs_3_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_3_io_inputs_0 = Alu_6_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_4_clock = clock;
  assign RegisterFiles_4_reset = reset;
  assign RegisterFiles_4_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_4_io_configuration = dispatchs_9_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_4_io_inputs_0 = Alu_7_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_5_clock = clock;
  assign RegisterFiles_5_reset = reset;
  assign RegisterFiles_5_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_5_io_configuration = dispatchs_6_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_5_io_inputs_0 = Alu_8_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_6_clock = clock;
  assign RegisterFiles_6_reset = reset;
  assign RegisterFiles_6_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_6_io_configuration = dispatchs_15_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_6_io_inputs_0 = Alu_9_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_7_clock = clock;
  assign RegisterFiles_7_reset = reset;
  assign RegisterFiles_7_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_7_io_configuration = dispatchs_18_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_7_io_inputs_0 = Alu_10_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_8_clock = clock;
  assign RegisterFiles_8_reset = reset;
  assign RegisterFiles_8_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_8_io_configuration = dispatchs_4_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_8_io_inputs_0 = Alu_11_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_9_clock = clock;
  assign RegisterFiles_9_reset = reset;
  assign RegisterFiles_9_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_9_io_configuration = dispatchs_10_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_9_io_inputs_0 = Alu_12_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_10_clock = clock;
  assign RegisterFiles_10_reset = reset;
  assign RegisterFiles_10_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_10_io_configuration = dispatchs_1_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_10_io_inputs_0 = Alu_13_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_11_clock = clock;
  assign RegisterFiles_11_reset = reset;
  assign RegisterFiles_11_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_11_io_configuration = dispatchs_20_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_11_io_inputs_0 = Alu_14_io_outs_0; // @[TopModule.scala 298:60]
  assign RegisterFiles_12_clock = clock;
  assign RegisterFiles_12_reset = reset;
  assign RegisterFiles_12_io_en = io_en; // @[TopModule.scala 148:14]
  assign RegisterFiles_12_io_configuration = dispatchs_8_io_outs_1; // @[TopModule.scala 249:22]
  assign RegisterFiles_12_io_inputs_0 = Alu_15_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_io_configuration = dispatchs_5_io_outs_0; // @[TopModule.scala 249:22]
  assign Multiplexer_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_1_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_1_io_configuration = dispatchs_5_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_1_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_1_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_1_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_1_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_2_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_2_io_configuration = dispatchs_5_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_2_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_2_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_2_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_2_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_3_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_3_io_configuration = dispatchs_5_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_3_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_3_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_3_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_3_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_4_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_4_io_configuration = dispatchs_5_io_outs_4; // @[TopModule.scala 249:22]
  assign Multiplexer_4_io_inputs_3 = io_inputs_3; // @[TopModule.scala 296:60]
  assign Multiplexer_4_io_inputs_2 = io_inputs_2; // @[TopModule.scala 296:60]
  assign Multiplexer_4_io_inputs_1 = io_inputs_1; // @[TopModule.scala 296:60]
  assign Multiplexer_4_io_inputs_0 = io_inputs_0; // @[TopModule.scala 296:60]
  assign Multiplexer_5_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_5_io_configuration = dispatchs_5_io_outs_5; // @[TopModule.scala 249:22]
  assign Multiplexer_5_io_inputs_3 = io_inputs_3; // @[TopModule.scala 296:60]
  assign Multiplexer_5_io_inputs_2 = io_inputs_2; // @[TopModule.scala 296:60]
  assign Multiplexer_5_io_inputs_1 = io_inputs_1; // @[TopModule.scala 296:60]
  assign Multiplexer_5_io_inputs_0 = io_inputs_0; // @[TopModule.scala 296:60]
  assign Multiplexer_6_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_6_io_configuration = dispatchs_5_io_outs_6; // @[TopModule.scala 249:22]
  assign Multiplexer_6_io_inputs_3 = io_inputs_3; // @[TopModule.scala 296:60]
  assign Multiplexer_6_io_inputs_2 = io_inputs_2; // @[TopModule.scala 296:60]
  assign Multiplexer_6_io_inputs_1 = io_inputs_1; // @[TopModule.scala 296:60]
  assign Multiplexer_6_io_inputs_0 = io_inputs_0; // @[TopModule.scala 296:60]
  assign Multiplexer_7_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_7_io_configuration = dispatchs_5_io_outs_7; // @[TopModule.scala 249:22]
  assign Multiplexer_7_io_inputs_3 = io_inputs_3; // @[TopModule.scala 296:60]
  assign Multiplexer_7_io_inputs_2 = io_inputs_2; // @[TopModule.scala 296:60]
  assign Multiplexer_7_io_inputs_1 = io_inputs_1; // @[TopModule.scala 296:60]
  assign Multiplexer_7_io_inputs_0 = io_inputs_0; // @[TopModule.scala 296:60]
  assign Multiplexer_8_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_8_io_configuration = dispatchs_2_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_8_io_inputs_7 = RegisterFiles_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_8_io_inputs_6 = ConstUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_8_io_inputs_5 = Multiplexer_4_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_8_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_8_io_inputs_3 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_8_io_inputs_2 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_8_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_8_io_inputs_0 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_9_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_9_io_configuration = dispatchs_2_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_9_io_inputs_6 = ConstUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_9_io_inputs_5 = Multiplexer_4_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_9_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_9_io_inputs_3 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_9_io_inputs_2 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_9_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_9_io_inputs_0 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_10_io_configuration = dispatchs_0_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_10_io_inputs_7 = RegisterFiles_io_outs_2; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_inputs_6 = ConstUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_inputs_5 = Multiplexer_5_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_inputs_3 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_inputs_2 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_inputs_1 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_10_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_11_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_11_io_configuration = dispatchs_0_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_11_io_inputs_6 = ConstUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_11_io_inputs_5 = Multiplexer_5_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_11_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_11_io_inputs_3 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_11_io_inputs_2 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_11_io_inputs_1 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_11_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_12_io_configuration = dispatchs_13_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_12_io_inputs_7 = RegisterFiles_io_outs_4; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_inputs_6 = ConstUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_inputs_5 = Multiplexer_6_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_inputs_3 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_inputs_2 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_inputs_1 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_12_io_inputs_0 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_13_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_13_io_configuration = dispatchs_13_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_13_io_inputs_6 = ConstUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_13_io_inputs_5 = Multiplexer_6_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_13_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_13_io_inputs_3 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_13_io_inputs_2 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_13_io_inputs_1 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_13_io_inputs_0 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_14_io_configuration = dispatchs_21_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_14_io_inputs_7 = RegisterFiles_io_outs_6; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_inputs_6 = ConstUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_inputs_5 = Multiplexer_7_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_inputs_3 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_inputs_2 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_inputs_1 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_14_io_inputs_0 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_15_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_15_io_configuration = dispatchs_21_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_15_io_inputs_6 = ConstUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_15_io_inputs_5 = Multiplexer_7_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_15_io_inputs_4 = LoadStoreUnit_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_15_io_inputs_3 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_15_io_inputs_2 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_15_io_inputs_1 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_15_io_inputs_0 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_16_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_16_io_configuration = dispatchs_12_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_16_io_inputs_6 = RegisterFiles_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_16_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_16_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_16_io_inputs_3 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_16_io_inputs_2 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_16_io_inputs_1 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_16_io_inputs_0 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_17_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_17_io_configuration = dispatchs_12_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_17_io_inputs_5 = ConstUnit_4_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_17_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_17_io_inputs_3 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_17_io_inputs_2 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_17_io_inputs_1 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_17_io_inputs_0 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_18_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_18_io_configuration = dispatchs_19_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_18_io_inputs_6 = RegisterFiles_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_18_io_inputs_5 = ConstUnit_5_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_18_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_18_io_inputs_3 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_18_io_inputs_2 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_18_io_inputs_1 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_18_io_inputs_0 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_19_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_19_io_configuration = dispatchs_19_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_19_io_inputs_5 = ConstUnit_5_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_19_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_19_io_inputs_3 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_19_io_inputs_2 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_19_io_inputs_1 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_19_io_inputs_0 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_20_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_20_io_configuration = dispatchs_3_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_20_io_inputs_6 = RegisterFiles_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_20_io_inputs_5 = ConstUnit_6_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_20_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_20_io_inputs_3 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_20_io_inputs_2 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_20_io_inputs_1 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_20_io_inputs_0 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_21_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_21_io_configuration = dispatchs_3_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_21_io_inputs_5 = ConstUnit_6_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_21_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_21_io_inputs_3 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_21_io_inputs_2 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_21_io_inputs_1 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_21_io_inputs_0 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_22_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_22_io_configuration = dispatchs_9_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_22_io_inputs_6 = RegisterFiles_4_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_22_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_22_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_22_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_22_io_inputs_2 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_22_io_inputs_1 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_22_io_inputs_0 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_23_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_23_io_configuration = dispatchs_9_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_23_io_inputs_5 = ConstUnit_7_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_23_io_inputs_4 = LoadStoreUnit_1_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_23_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_23_io_inputs_2 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_23_io_inputs_1 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_23_io_inputs_0 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_24_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_24_io_configuration = dispatchs_6_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_24_io_inputs_6 = RegisterFiles_5_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_24_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_24_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_24_io_inputs_3 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_24_io_inputs_2 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_24_io_inputs_1 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_24_io_inputs_0 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_25_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_25_io_configuration = dispatchs_6_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_25_io_inputs_5 = ConstUnit_8_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_25_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_25_io_inputs_3 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_25_io_inputs_2 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_25_io_inputs_1 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_25_io_inputs_0 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_26_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_26_io_configuration = dispatchs_15_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_26_io_inputs_6 = RegisterFiles_6_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_26_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_26_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_26_io_inputs_3 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_26_io_inputs_2 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_26_io_inputs_1 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_26_io_inputs_0 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_27_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_27_io_configuration = dispatchs_15_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_27_io_inputs_5 = ConstUnit_9_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_27_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_27_io_inputs_3 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_27_io_inputs_2 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_27_io_inputs_1 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_27_io_inputs_0 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_28_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_28_io_configuration = dispatchs_18_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_28_io_inputs_6 = RegisterFiles_7_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_28_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_28_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_28_io_inputs_3 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_28_io_inputs_2 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_28_io_inputs_1 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_28_io_inputs_0 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_29_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_29_io_configuration = dispatchs_18_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_29_io_inputs_5 = ConstUnit_10_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_29_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_29_io_inputs_3 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_29_io_inputs_2 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_29_io_inputs_1 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_29_io_inputs_0 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_30_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_30_io_configuration = dispatchs_4_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_30_io_inputs_6 = RegisterFiles_8_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_30_io_inputs_5 = ConstUnit_11_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_30_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_30_io_inputs_3 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_30_io_inputs_2 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_30_io_inputs_1 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_30_io_inputs_0 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_31_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_31_io_configuration = dispatchs_4_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_31_io_inputs_5 = ConstUnit_11_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_31_io_inputs_4 = LoadStoreUnit_2_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_31_io_inputs_3 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_31_io_inputs_2 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_31_io_inputs_1 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_31_io_inputs_0 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_32_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_32_io_configuration = dispatchs_10_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_32_io_inputs_6 = RegisterFiles_9_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_32_io_inputs_5 = ConstUnit_12_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_32_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_32_io_inputs_3 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_32_io_inputs_2 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_32_io_inputs_1 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_32_io_inputs_0 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_33_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_33_io_configuration = dispatchs_10_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_33_io_inputs_5 = ConstUnit_12_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_33_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_33_io_inputs_3 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_33_io_inputs_2 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_33_io_inputs_1 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_33_io_inputs_0 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_34_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_34_io_configuration = dispatchs_1_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_34_io_inputs_6 = RegisterFiles_10_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_34_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_34_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_34_io_inputs_3 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_34_io_inputs_2 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_34_io_inputs_1 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_34_io_inputs_0 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_35_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_35_io_configuration = dispatchs_1_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_35_io_inputs_5 = ConstUnit_13_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_35_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_35_io_inputs_3 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_35_io_inputs_2 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_35_io_inputs_1 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_35_io_inputs_0 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_36_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_36_io_configuration = dispatchs_20_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_36_io_inputs_6 = RegisterFiles_11_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_36_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_36_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_36_io_inputs_3 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_36_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_36_io_inputs_1 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_36_io_inputs_0 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_37_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_37_io_configuration = dispatchs_20_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_37_io_inputs_5 = ConstUnit_14_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_37_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_37_io_inputs_3 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_37_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_37_io_inputs_1 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_37_io_inputs_0 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_38_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_38_io_configuration = dispatchs_8_io_outs_2; // @[TopModule.scala 249:22]
  assign Multiplexer_38_io_inputs_6 = RegisterFiles_12_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_38_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_38_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_38_io_inputs_3 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_38_io_inputs_2 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_38_io_inputs_1 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_38_io_inputs_0 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_39_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_39_io_configuration = dispatchs_8_io_outs_3; // @[TopModule.scala 249:22]
  assign Multiplexer_39_io_inputs_5 = ConstUnit_15_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_39_io_inputs_4 = LoadStoreUnit_3_io_outs_0; // @[TopModule.scala 298:60]
  assign Multiplexer_39_io_inputs_3 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_39_io_inputs_2 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_39_io_inputs_1 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_39_io_inputs_0 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_40_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_40_io_configuration = dispatchs_7_io_outs_0; // @[TopModule.scala 249:22]
  assign Multiplexer_40_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_40_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_40_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_40_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_41_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_41_io_configuration = dispatchs_7_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_41_io_inputs_3 = RegisterFiles_io_outs_7; // @[TopModule.scala 298:60]
  assign Multiplexer_41_io_inputs_2 = RegisterFiles_io_outs_5; // @[TopModule.scala 298:60]
  assign Multiplexer_41_io_inputs_1 = RegisterFiles_io_outs_3; // @[TopModule.scala 298:60]
  assign Multiplexer_41_io_inputs_0 = RegisterFiles_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_42_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_42_io_configuration = dispatchs_14_io_outs_0; // @[TopModule.scala 249:22]
  assign Multiplexer_42_io_inputs_3 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_42_io_inputs_2 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_42_io_inputs_1 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_42_io_inputs_0 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_43_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_43_io_configuration = dispatchs_14_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_43_io_inputs_3 = RegisterFiles_4_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_43_io_inputs_2 = RegisterFiles_3_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_43_io_inputs_1 = RegisterFiles_2_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_43_io_inputs_0 = RegisterFiles_1_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_44_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_44_io_configuration = dispatchs_17_io_outs_0; // @[TopModule.scala 249:22]
  assign Multiplexer_44_io_inputs_3 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_44_io_inputs_2 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_44_io_inputs_1 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_44_io_inputs_0 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_45_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_45_io_configuration = dispatchs_17_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_45_io_inputs_3 = RegisterFiles_8_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_45_io_inputs_2 = RegisterFiles_7_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_45_io_inputs_1 = RegisterFiles_6_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_45_io_inputs_0 = RegisterFiles_5_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_46_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_46_io_configuration = dispatchs_11_io_outs_0; // @[TopModule.scala 249:22]
  assign Multiplexer_46_io_inputs_3 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_46_io_inputs_2 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_46_io_inputs_1 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_46_io_inputs_0 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_47_io_en = io_en; // @[TopModule.scala 157:15]
  assign Multiplexer_47_io_configuration = dispatchs_11_io_outs_1; // @[TopModule.scala 249:22]
  assign Multiplexer_47_io_inputs_3 = RegisterFiles_12_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_47_io_inputs_2 = RegisterFiles_11_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_47_io_inputs_1 = RegisterFiles_10_io_outs_1; // @[TopModule.scala 298:60]
  assign Multiplexer_47_io_inputs_0 = RegisterFiles_9_io_outs_1; // @[TopModule.scala 298:60]
  assign ConstUnit_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_io_configuration = dispatchs_2_io_outs_3; // @[TopModule.scala 249:22]
  assign ConstUnit_1_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_1_io_configuration = dispatchs_0_io_outs_3; // @[TopModule.scala 249:22]
  assign ConstUnit_2_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_2_io_configuration = dispatchs_13_io_outs_3; // @[TopModule.scala 249:22]
  assign ConstUnit_3_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_3_io_configuration = dispatchs_21_io_outs_3; // @[TopModule.scala 249:22]
  assign ConstUnit_4_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_4_io_configuration = dispatchs_12_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_5_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_5_io_configuration = dispatchs_19_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_6_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_6_io_configuration = dispatchs_3_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_7_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_7_io_configuration = dispatchs_9_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_8_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_8_io_configuration = dispatchs_6_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_9_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_9_io_configuration = dispatchs_15_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_10_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_10_io_configuration = dispatchs_18_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_11_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_11_io_configuration = dispatchs_4_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_12_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_12_io_configuration = dispatchs_10_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_13_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_13_io_configuration = dispatchs_1_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_14_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_14_io_configuration = dispatchs_20_io_outs_4; // @[TopModule.scala 249:22]
  assign ConstUnit_15_io_en = io_en; // @[TopModule.scala 165:17]
  assign ConstUnit_15_io_configuration = dispatchs_8_io_outs_4; // @[TopModule.scala 249:22]
  assign LoadStoreUnit_clock = clock;
  assign LoadStoreUnit_reset = reset;
  assign LoadStoreUnit_io_configuration = dispatchs_7_io_outs_2; // @[TopModule.scala 249:22]
  assign LoadStoreUnit_io_en = MultiIIScheduleController_16_io_valid; // @[TopModule.scala 194:15]
  assign LoadStoreUnit_io_skewing = MultiIIScheduleController_16_io_skewing; // @[TopModule.scala 195:20]
  assign LoadStoreUnit_io_streamIn_valid = io_streamInLSU_0_valid; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_io_streamIn_bits = io_streamInLSU_0_bits; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_io_len = io_lenLSU_0; // @[TopModule.scala 179:16]
  assign LoadStoreUnit_io_streamOut_ready = io_streamOutLSU_0_ready; // @[TopModule.scala 185:22]
  assign LoadStoreUnit_io_base = io_baseLSU_0; // @[TopModule.scala 178:17]
  assign LoadStoreUnit_io_start = io_startLSU_0; // @[TopModule.scala 180:18]
  assign LoadStoreUnit_io_enqEn = io_enqEnLSU_0; // @[TopModule.scala 182:18]
  assign LoadStoreUnit_io_deqEn = io_deqEnLSU_0; // @[TopModule.scala 183:18]
  assign LoadStoreUnit_io_inputs_1 = Multiplexer_41_io_outs_0; // @[TopModule.scala 298:60]
  assign LoadStoreUnit_io_inputs_0 = Multiplexer_40_io_outs_0[7:0]; // @[TopModule.scala 298:60]
  assign LoadStoreUnit_1_clock = clock;
  assign LoadStoreUnit_1_reset = reset;
  assign LoadStoreUnit_1_io_configuration = dispatchs_14_io_outs_2; // @[TopModule.scala 249:22]
  assign LoadStoreUnit_1_io_en = MultiIIScheduleController_17_io_valid; // @[TopModule.scala 194:15]
  assign LoadStoreUnit_1_io_skewing = MultiIIScheduleController_17_io_skewing; // @[TopModule.scala 195:20]
  assign LoadStoreUnit_1_io_streamIn_valid = io_streamInLSU_1_valid; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_1_io_streamIn_bits = io_streamInLSU_1_bits; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_1_io_len = io_lenLSU_1; // @[TopModule.scala 179:16]
  assign LoadStoreUnit_1_io_streamOut_ready = io_streamOutLSU_1_ready; // @[TopModule.scala 185:22]
  assign LoadStoreUnit_1_io_base = io_baseLSU_1; // @[TopModule.scala 178:17]
  assign LoadStoreUnit_1_io_start = io_startLSU_1; // @[TopModule.scala 180:18]
  assign LoadStoreUnit_1_io_enqEn = io_enqEnLSU_1; // @[TopModule.scala 182:18]
  assign LoadStoreUnit_1_io_deqEn = io_deqEnLSU_1; // @[TopModule.scala 183:18]
  assign LoadStoreUnit_1_io_inputs_1 = Multiplexer_43_io_outs_0; // @[TopModule.scala 298:60]
  assign LoadStoreUnit_1_io_inputs_0 = Multiplexer_42_io_outs_0[7:0]; // @[TopModule.scala 298:60]
  assign LoadStoreUnit_2_clock = clock;
  assign LoadStoreUnit_2_reset = reset;
  assign LoadStoreUnit_2_io_configuration = dispatchs_17_io_outs_2; // @[TopModule.scala 249:22]
  assign LoadStoreUnit_2_io_en = MultiIIScheduleController_18_io_valid; // @[TopModule.scala 194:15]
  assign LoadStoreUnit_2_io_skewing = MultiIIScheduleController_18_io_skewing; // @[TopModule.scala 195:20]
  assign LoadStoreUnit_2_io_streamIn_valid = io_streamInLSU_2_valid; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_2_io_streamIn_bits = io_streamInLSU_2_bits; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_2_io_len = io_lenLSU_2; // @[TopModule.scala 179:16]
  assign LoadStoreUnit_2_io_streamOut_ready = io_streamOutLSU_2_ready; // @[TopModule.scala 185:22]
  assign LoadStoreUnit_2_io_base = io_baseLSU_2; // @[TopModule.scala 178:17]
  assign LoadStoreUnit_2_io_start = io_startLSU_2; // @[TopModule.scala 180:18]
  assign LoadStoreUnit_2_io_enqEn = io_enqEnLSU_2; // @[TopModule.scala 182:18]
  assign LoadStoreUnit_2_io_deqEn = io_deqEnLSU_2; // @[TopModule.scala 183:18]
  assign LoadStoreUnit_2_io_inputs_1 = Multiplexer_45_io_outs_0; // @[TopModule.scala 298:60]
  assign LoadStoreUnit_2_io_inputs_0 = Multiplexer_44_io_outs_0[7:0]; // @[TopModule.scala 298:60]
  assign LoadStoreUnit_3_clock = clock;
  assign LoadStoreUnit_3_reset = reset;
  assign LoadStoreUnit_3_io_configuration = dispatchs_11_io_outs_2; // @[TopModule.scala 249:22]
  assign LoadStoreUnit_3_io_en = MultiIIScheduleController_19_io_valid; // @[TopModule.scala 194:15]
  assign LoadStoreUnit_3_io_skewing = MultiIIScheduleController_19_io_skewing; // @[TopModule.scala 195:20]
  assign LoadStoreUnit_3_io_streamIn_valid = io_streamInLSU_3_valid; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_3_io_streamIn_bits = io_streamInLSU_3_bits; // @[TopModule.scala 184:21]
  assign LoadStoreUnit_3_io_len = io_lenLSU_3; // @[TopModule.scala 179:16]
  assign LoadStoreUnit_3_io_streamOut_ready = io_streamOutLSU_3_ready; // @[TopModule.scala 185:22]
  assign LoadStoreUnit_3_io_base = io_baseLSU_3; // @[TopModule.scala 178:17]
  assign LoadStoreUnit_3_io_start = io_startLSU_3; // @[TopModule.scala 180:18]
  assign LoadStoreUnit_3_io_enqEn = io_enqEnLSU_3; // @[TopModule.scala 182:18]
  assign LoadStoreUnit_3_io_deqEn = io_deqEnLSU_3; // @[TopModule.scala 183:18]
  assign LoadStoreUnit_3_io_inputs_1 = Multiplexer_47_io_outs_0; // @[TopModule.scala 298:60]
  assign LoadStoreUnit_3_io_inputs_0 = Multiplexer_46_io_outs_0[7:0]; // @[TopModule.scala 298:60]
  assign MultiIIScheduleController_16_clock = clock;
  assign MultiIIScheduleController_16_reset = reset;
  assign MultiIIScheduleController_16_io_en = io_en; // @[TopModule.scala 189:36]
  assign MultiIIScheduleController_16_io_schedules_0 = 9'h0; // @[TopModule.scala 192:48]
  assign MultiIIScheduleController_16_io_II = io_II; // @[TopModule.scala 190:36]
  assign MultiIIScheduleController_17_clock = clock;
  assign MultiIIScheduleController_17_reset = reset;
  assign MultiIIScheduleController_17_io_en = io_en; // @[TopModule.scala 189:36]
  assign MultiIIScheduleController_17_io_schedules_0 = 9'h0; // @[TopModule.scala 192:48]
  assign MultiIIScheduleController_17_io_II = io_II; // @[TopModule.scala 190:36]
  assign MultiIIScheduleController_18_clock = clock;
  assign MultiIIScheduleController_18_reset = reset;
  assign MultiIIScheduleController_18_io_en = io_en; // @[TopModule.scala 189:36]
  assign MultiIIScheduleController_18_io_schedules_0 = scheduleDispatch_io_outs_144; // @[TopModule.scala 192:48]
  assign MultiIIScheduleController_18_io_II = io_II; // @[TopModule.scala 190:36]
  assign MultiIIScheduleController_19_clock = clock;
  assign MultiIIScheduleController_19_reset = reset;
  assign MultiIIScheduleController_19_io_en = io_en; // @[TopModule.scala 189:36]
  assign MultiIIScheduleController_19_io_schedules_0 = 9'h0; // @[TopModule.scala 192:48]
  assign MultiIIScheduleController_19_io_II = io_II; // @[TopModule.scala 190:36]
  assign configController_clock = clock;
  assign configController_reset = reset;
  assign configController_io_en = io_en; // @[TopModule.scala 220:26]
  assign configController_io_II = io_II; // @[TopModule.scala 221:26]
  assign dispatchs_0_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_0_io_configuration = topDispatch_io_outs_0; // @[TopModule.scala 261:35]
  assign dispatchs_1_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_1_io_configuration = topDispatch_io_outs_1; // @[TopModule.scala 261:35]
  assign dispatchs_2_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_2_io_configuration = topDispatch_io_outs_2; // @[TopModule.scala 261:35]
  assign dispatchs_3_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_3_io_configuration = topDispatch_io_outs_3; // @[TopModule.scala 261:35]
  assign dispatchs_4_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_4_io_configuration = topDispatch_io_outs_4; // @[TopModule.scala 261:35]
  assign dispatchs_5_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_5_io_configuration = topDispatch_io_outs_5; // @[TopModule.scala 261:35]
  assign dispatchs_6_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_6_io_configuration = topDispatch_io_outs_6; // @[TopModule.scala 261:35]
  assign dispatchs_7_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_7_io_configuration = topDispatch_io_outs_7; // @[TopModule.scala 261:35]
  assign dispatchs_8_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_8_io_configuration = topDispatch_io_outs_8; // @[TopModule.scala 261:35]
  assign dispatchs_9_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_9_io_configuration = topDispatch_io_outs_9; // @[TopModule.scala 261:35]
  assign dispatchs_10_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_10_io_configuration = topDispatch_io_outs_10; // @[TopModule.scala 261:35]
  assign dispatchs_11_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_11_io_configuration = topDispatch_io_outs_11; // @[TopModule.scala 261:35]
  assign dispatchs_12_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_12_io_configuration = topDispatch_io_outs_12; // @[TopModule.scala 261:35]
  assign dispatchs_13_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_13_io_configuration = topDispatch_io_outs_13; // @[TopModule.scala 261:35]
  assign dispatchs_14_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_14_io_configuration = topDispatch_io_outs_14; // @[TopModule.scala 261:35]
  assign dispatchs_15_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_15_io_configuration = topDispatch_io_outs_15; // @[TopModule.scala 261:35]
  assign dispatchs_16_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_16_io_configuration = topDispatch_io_outs_16; // @[TopModule.scala 261:35]
  assign dispatchs_17_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_17_io_configuration = topDispatch_io_outs_17; // @[TopModule.scala 261:35]
  assign dispatchs_18_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_18_io_configuration = topDispatch_io_outs_18; // @[TopModule.scala 261:35]
  assign dispatchs_19_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_19_io_configuration = topDispatch_io_outs_19; // @[TopModule.scala 261:35]
  assign dispatchs_20_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_20_io_configuration = topDispatch_io_outs_20; // @[TopModule.scala 261:35]
  assign dispatchs_21_io_en = io_en; // @[TopModule.scala 247:20]
  assign dispatchs_21_io_configuration = topDispatch_io_outs_21; // @[TopModule.scala 261:35]
  assign topDispatch_io_en = io_en; // @[TopModule.scala 256:21]
  assign topDispatch_io_configuration = configController_io_outConfig; // @[TopModule.scala 259:32]
endmodule
module TopModuleWrapper(
  input         clock,
  input         reset,
  output        io_streamInLSU_ready,
  input         io_streamInLSU_valid,
  input  [31:0] io_streamInLSU_bits,
  input         io_streamOutLSU_ready,
  output        io_streamOutLSU_valid,
  output [31:0] io_streamOutLSU_bits,
  input  [7:0]  io_baseLSU,
  input  [7:0]  io_lenLSU,
  input         io_startLSU,
  input         io_enqEnLSU,
  input         io_deqEnLSU,
  output        io_idleLSU,
  input  [1:0]  io_LSUnitID,
  input         io_en,
  input  [2:0]  io_II,
  input  [31:0] io_inputs_3,
  input  [31:0] io_inputs_2,
  input  [31:0] io_inputs_1,
  input  [31:0] io_inputs_0,
  output [31:0] io_outs_3,
  output [31:0] io_outs_2,
  output [31:0] io_outs_1,
  output [31:0] io_outs_0
);
  wire  topModule_clock; // @[TopModule.scala 310:25]
  wire  topModule_reset; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_3_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_3_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamInLSU_3_bits; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_2_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_2_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamInLSU_2_bits; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_1_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_1_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamInLSU_1_bits; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_0_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamInLSU_0_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamInLSU_0_bits; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_3_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_3_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamOutLSU_3_bits; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_2_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_2_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamOutLSU_2_bits; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_1_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_1_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamOutLSU_1_bits; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_0_ready; // @[TopModule.scala 310:25]
  wire  topModule_io_streamOutLSU_0_valid; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_streamOutLSU_0_bits; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_baseLSU_0; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_baseLSU_1; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_baseLSU_2; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_baseLSU_3; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_lenLSU_0; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_lenLSU_1; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_lenLSU_2; // @[TopModule.scala 310:25]
  wire [7:0] topModule_io_lenLSU_3; // @[TopModule.scala 310:25]
  wire  topModule_io_startLSU_0; // @[TopModule.scala 310:25]
  wire  topModule_io_startLSU_1; // @[TopModule.scala 310:25]
  wire  topModule_io_startLSU_2; // @[TopModule.scala 310:25]
  wire  topModule_io_startLSU_3; // @[TopModule.scala 310:25]
  wire  topModule_io_enqEnLSU_0; // @[TopModule.scala 310:25]
  wire  topModule_io_enqEnLSU_1; // @[TopModule.scala 310:25]
  wire  topModule_io_enqEnLSU_2; // @[TopModule.scala 310:25]
  wire  topModule_io_enqEnLSU_3; // @[TopModule.scala 310:25]
  wire  topModule_io_deqEnLSU_0; // @[TopModule.scala 310:25]
  wire  topModule_io_deqEnLSU_1; // @[TopModule.scala 310:25]
  wire  topModule_io_deqEnLSU_2; // @[TopModule.scala 310:25]
  wire  topModule_io_deqEnLSU_3; // @[TopModule.scala 310:25]
  wire  topModule_io_idleLSU_0; // @[TopModule.scala 310:25]
  wire  topModule_io_idleLSU_1; // @[TopModule.scala 310:25]
  wire  topModule_io_idleLSU_2; // @[TopModule.scala 310:25]
  wire  topModule_io_idleLSU_3; // @[TopModule.scala 310:25]
  wire  topModule_io_en; // @[TopModule.scala 310:25]
  wire [2:0] topModule_io_II; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_inputs_3; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_inputs_2; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_inputs_1; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_inputs_0; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_outs_3; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_outs_2; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_outs_1; // @[TopModule.scala 310:25]
  wire [31:0] topModule_io_outs_0; // @[TopModule.scala 310:25]
  wire  _T; // @[TopModule.scala 358:20]
  wire  _T_1; // @[TopModule.scala 360:26]
  wire  _T_2; // @[TopModule.scala 362:26]
  wire [31:0] _GEN_5; // @[TopModule.scala 362:34]
  wire  _GEN_6; // @[TopModule.scala 362:34]
  wire [31:0] _GEN_8; // @[TopModule.scala 362:34]
  wire  _GEN_9; // @[TopModule.scala 362:34]
  wire  _GEN_10; // @[TopModule.scala 362:34]
  wire  _GEN_18; // @[TopModule.scala 362:34]
  wire [31:0] _GEN_19; // @[TopModule.scala 362:34]
  wire [31:0] _GEN_25; // @[TopModule.scala 360:34]
  wire  _GEN_26; // @[TopModule.scala 360:34]
  wire [31:0] _GEN_28; // @[TopModule.scala 360:34]
  wire  _GEN_29; // @[TopModule.scala 360:34]
  wire  _GEN_30; // @[TopModule.scala 360:34]
  wire  _GEN_38; // @[TopModule.scala 360:34]
  wire [31:0] _GEN_39; // @[TopModule.scala 360:34]
  wire  _GEN_46; // @[TopModule.scala 360:34]
  wire [31:0] _GEN_47; // @[TopModule.scala 360:34]
  wire  _GEN_83; // @[TopModule.scala 368:37]
  wire  _GEN_84; // @[TopModule.scala 368:37]
  wire  _GEN_85; // @[TopModule.scala 368:37]
  TopModule topModule ( // @[TopModule.scala 310:25]
    .clock(topModule_clock),
    .reset(topModule_reset),
    .io_streamInLSU_3_ready(topModule_io_streamInLSU_3_ready),
    .io_streamInLSU_3_valid(topModule_io_streamInLSU_3_valid),
    .io_streamInLSU_3_bits(topModule_io_streamInLSU_3_bits),
    .io_streamInLSU_2_ready(topModule_io_streamInLSU_2_ready),
    .io_streamInLSU_2_valid(topModule_io_streamInLSU_2_valid),
    .io_streamInLSU_2_bits(topModule_io_streamInLSU_2_bits),
    .io_streamInLSU_1_ready(topModule_io_streamInLSU_1_ready),
    .io_streamInLSU_1_valid(topModule_io_streamInLSU_1_valid),
    .io_streamInLSU_1_bits(topModule_io_streamInLSU_1_bits),
    .io_streamInLSU_0_ready(topModule_io_streamInLSU_0_ready),
    .io_streamInLSU_0_valid(topModule_io_streamInLSU_0_valid),
    .io_streamInLSU_0_bits(topModule_io_streamInLSU_0_bits),
    .io_streamOutLSU_3_ready(topModule_io_streamOutLSU_3_ready),
    .io_streamOutLSU_3_valid(topModule_io_streamOutLSU_3_valid),
    .io_streamOutLSU_3_bits(topModule_io_streamOutLSU_3_bits),
    .io_streamOutLSU_2_ready(topModule_io_streamOutLSU_2_ready),
    .io_streamOutLSU_2_valid(topModule_io_streamOutLSU_2_valid),
    .io_streamOutLSU_2_bits(topModule_io_streamOutLSU_2_bits),
    .io_streamOutLSU_1_ready(topModule_io_streamOutLSU_1_ready),
    .io_streamOutLSU_1_valid(topModule_io_streamOutLSU_1_valid),
    .io_streamOutLSU_1_bits(topModule_io_streamOutLSU_1_bits),
    .io_streamOutLSU_0_ready(topModule_io_streamOutLSU_0_ready),
    .io_streamOutLSU_0_valid(topModule_io_streamOutLSU_0_valid),
    .io_streamOutLSU_0_bits(topModule_io_streamOutLSU_0_bits),
    .io_baseLSU_0(topModule_io_baseLSU_0),
    .io_baseLSU_1(topModule_io_baseLSU_1),
    .io_baseLSU_2(topModule_io_baseLSU_2),
    .io_baseLSU_3(topModule_io_baseLSU_3),
    .io_lenLSU_0(topModule_io_lenLSU_0),
    .io_lenLSU_1(topModule_io_lenLSU_1),
    .io_lenLSU_2(topModule_io_lenLSU_2),
    .io_lenLSU_3(topModule_io_lenLSU_3),
    .io_startLSU_0(topModule_io_startLSU_0),
    .io_startLSU_1(topModule_io_startLSU_1),
    .io_startLSU_2(topModule_io_startLSU_2),
    .io_startLSU_3(topModule_io_startLSU_3),
    .io_enqEnLSU_0(topModule_io_enqEnLSU_0),
    .io_enqEnLSU_1(topModule_io_enqEnLSU_1),
    .io_enqEnLSU_2(topModule_io_enqEnLSU_2),
    .io_enqEnLSU_3(topModule_io_enqEnLSU_3),
    .io_deqEnLSU_0(topModule_io_deqEnLSU_0),
    .io_deqEnLSU_1(topModule_io_deqEnLSU_1),
    .io_deqEnLSU_2(topModule_io_deqEnLSU_2),
    .io_deqEnLSU_3(topModule_io_deqEnLSU_3),
    .io_idleLSU_0(topModule_io_idleLSU_0),
    .io_idleLSU_1(topModule_io_idleLSU_1),
    .io_idleLSU_2(topModule_io_idleLSU_2),
    .io_idleLSU_3(topModule_io_idleLSU_3),
    .io_en(topModule_io_en),
    .io_II(topModule_io_II),
    .io_inputs_3(topModule_io_inputs_3),
    .io_inputs_2(topModule_io_inputs_2),
    .io_inputs_1(topModule_io_inputs_1),
    .io_inputs_0(topModule_io_inputs_0),
    .io_outs_3(topModule_io_outs_3),
    .io_outs_2(topModule_io_outs_2),
    .io_outs_1(topModule_io_outs_1),
    .io_outs_0(topModule_io_outs_0)
  );
  assign _T = io_LSUnitID == 2'h0; // @[TopModule.scala 358:20]
  assign _T_1 = io_LSUnitID == 2'h1; // @[TopModule.scala 360:26]
  assign _T_2 = io_LSUnitID == 2'h2; // @[TopModule.scala 362:26]
  assign _GEN_5 = _T_2 ? topModule_io_streamOutLSU_2_bits : topModule_io_streamOutLSU_3_bits; // @[TopModule.scala 362:34]
  assign _GEN_6 = _T_2 ? topModule_io_streamOutLSU_2_valid : topModule_io_streamOutLSU_3_valid; // @[TopModule.scala 362:34]
  assign _GEN_8 = _T_2 ? io_streamInLSU_bits : 32'h0; // @[TopModule.scala 362:34]
  assign _GEN_9 = _T_2 & io_streamInLSU_valid; // @[TopModule.scala 362:34]
  assign _GEN_10 = _T_2 ? topModule_io_streamInLSU_2_ready : topModule_io_streamInLSU_3_ready; // @[TopModule.scala 362:34]
  assign _GEN_18 = _T_2 ? 1'h0 : io_streamInLSU_valid; // @[TopModule.scala 362:34]
  assign _GEN_19 = _T_2 ? 32'h0 : io_streamInLSU_bits; // @[TopModule.scala 362:34]
  assign _GEN_25 = _T_1 ? topModule_io_streamOutLSU_1_bits : _GEN_5; // @[TopModule.scala 360:34]
  assign _GEN_26 = _T_1 ? topModule_io_streamOutLSU_1_valid : _GEN_6; // @[TopModule.scala 360:34]
  assign _GEN_28 = _T_1 ? io_streamInLSU_bits : 32'h0; // @[TopModule.scala 360:34]
  assign _GEN_29 = _T_1 & io_streamInLSU_valid; // @[TopModule.scala 360:34]
  assign _GEN_30 = _T_1 ? topModule_io_streamInLSU_1_ready : _GEN_10; // @[TopModule.scala 360:34]
  assign _GEN_38 = _T_1 ? 1'h0 : _GEN_9; // @[TopModule.scala 360:34]
  assign _GEN_39 = _T_1 ? 32'h0 : _GEN_8; // @[TopModule.scala 360:34]
  assign _GEN_46 = _T_1 ? 1'h0 : _GEN_18; // @[TopModule.scala 360:34]
  assign _GEN_47 = _T_1 ? 32'h0 : _GEN_19; // @[TopModule.scala 360:34]
  assign _GEN_83 = topModule_io_idleLSU_0; // @[TopModule.scala 368:37]
  assign _GEN_84 = 2'h1 == io_LSUnitID ? topModule_io_idleLSU_1 : _GEN_83; // @[TopModule.scala 368:37]
  assign _GEN_85 = 2'h2 == io_LSUnitID ? topModule_io_idleLSU_2 : _GEN_84; // @[TopModule.scala 368:37]
  assign io_streamInLSU_ready = _T ? topModule_io_streamInLSU_0_ready : _GEN_30; // @[TopModule.scala 343:33 TopModule.scala 343:33 TopModule.scala 343:33 TopModule.scala 343:33]
  assign io_streamOutLSU_valid = _T ? topModule_io_streamOutLSU_0_valid : _GEN_26; // @[TopModule.scala 342:34 TopModule.scala 342:34 TopModule.scala 342:34 TopModule.scala 342:34]
  assign io_streamOutLSU_bits = _T ? topModule_io_streamOutLSU_0_bits : _GEN_25; // @[TopModule.scala 342:34 TopModule.scala 342:34 TopModule.scala 342:34 TopModule.scala 342:34]
  assign io_idleLSU = 2'h3 == io_LSUnitID ? topModule_io_idleLSU_3 : _GEN_85; // @[TopModule.scala 368:37]
  assign io_outs_3 = topModule_io_outs_3; // @[TopModule.scala 371:21]
  assign io_outs_2 = topModule_io_outs_2; // @[TopModule.scala 371:21]
  assign io_outs_1 = topModule_io_outs_1; // @[TopModule.scala 371:21]
  assign io_outs_0 = topModule_io_outs_0; // @[TopModule.scala 371:21]
  assign topModule_clock = clock;
  assign topModule_reset = reset;
  assign topModule_io_streamInLSU_3_valid = _T ? 1'h0 : _GEN_46; // @[TopModule.scala 352:43 TopModule.scala 352:43 TopModule.scala 352:43 TopModule.scala 343:33]
  assign topModule_io_streamInLSU_3_bits = _T ? 32'h0 : _GEN_47; // @[TopModule.scala 353:42 TopModule.scala 353:42 TopModule.scala 353:42 TopModule.scala 343:33]
  assign topModule_io_streamInLSU_2_valid = _T ? 1'h0 : _GEN_38; // @[TopModule.scala 352:43 TopModule.scala 352:43 TopModule.scala 343:33 TopModule.scala 352:43]
  assign topModule_io_streamInLSU_2_bits = _T ? 32'h0 : _GEN_39; // @[TopModule.scala 353:42 TopModule.scala 353:42 TopModule.scala 343:33 TopModule.scala 353:42]
  assign topModule_io_streamInLSU_1_valid = _T ? 1'h0 : _GEN_29; // @[TopModule.scala 352:43 TopModule.scala 343:33 TopModule.scala 352:43 TopModule.scala 352:43]
  assign topModule_io_streamInLSU_1_bits = _T ? 32'h0 : _GEN_28; // @[TopModule.scala 353:42 TopModule.scala 343:33 TopModule.scala 353:42 TopModule.scala 353:42]
  assign topModule_io_streamInLSU_0_valid = _T & io_streamInLSU_valid; // @[TopModule.scala 343:33 TopModule.scala 352:43 TopModule.scala 352:43 TopModule.scala 352:43]
  assign topModule_io_streamInLSU_0_bits = _T ? io_streamInLSU_bits : 32'h0; // @[TopModule.scala 343:33 TopModule.scala 353:42 TopModule.scala 353:42 TopModule.scala 353:42]
  assign topModule_io_streamOutLSU_3_ready = io_streamOutLSU_ready; // @[TopModule.scala 342:34]
  assign topModule_io_streamOutLSU_2_ready = io_streamOutLSU_ready; // @[TopModule.scala 342:34]
  assign topModule_io_streamOutLSU_1_ready = io_streamOutLSU_ready; // @[TopModule.scala 342:34]
  assign topModule_io_streamOutLSU_0_ready = io_streamOutLSU_ready; // @[TopModule.scala 342:34]
  assign topModule_io_baseLSU_0 = io_baseLSU; // @[TopModule.scala 337:31]
  assign topModule_io_baseLSU_1 = io_baseLSU; // @[TopModule.scala 337:31]
  assign topModule_io_baseLSU_2 = io_baseLSU; // @[TopModule.scala 337:31]
  assign topModule_io_baseLSU_3 = io_baseLSU; // @[TopModule.scala 337:31]
  assign topModule_io_lenLSU_0 = io_lenLSU; // @[TopModule.scala 338:30]
  assign topModule_io_lenLSU_1 = io_lenLSU; // @[TopModule.scala 338:30]
  assign topModule_io_lenLSU_2 = io_lenLSU; // @[TopModule.scala 338:30]
  assign topModule_io_lenLSU_3 = io_lenLSU; // @[TopModule.scala 338:30]
  assign topModule_io_startLSU_0 = io_startLSU; // @[TopModule.scala 339:32]
  assign topModule_io_startLSU_1 = io_startLSU; // @[TopModule.scala 339:32]
  assign topModule_io_startLSU_2 = io_startLSU; // @[TopModule.scala 339:32]
  assign topModule_io_startLSU_3 = io_startLSU; // @[TopModule.scala 339:32]
  assign topModule_io_enqEnLSU_0 = io_enqEnLSU; // @[TopModule.scala 340:32]
  assign topModule_io_enqEnLSU_1 = io_enqEnLSU; // @[TopModule.scala 340:32]
  assign topModule_io_enqEnLSU_2 = io_enqEnLSU; // @[TopModule.scala 340:32]
  assign topModule_io_enqEnLSU_3 = io_enqEnLSU; // @[TopModule.scala 340:32]
  assign topModule_io_deqEnLSU_0 = io_deqEnLSU; // @[TopModule.scala 341:32]
  assign topModule_io_deqEnLSU_1 = io_deqEnLSU; // @[TopModule.scala 341:32]
  assign topModule_io_deqEnLSU_2 = io_deqEnLSU; // @[TopModule.scala 341:32]
  assign topModule_io_deqEnLSU_3 = io_deqEnLSU; // @[TopModule.scala 341:32]
  assign topModule_io_en = io_en; // @[TopModule.scala 333:19]
  assign topModule_io_II = io_II; // @[TopModule.scala 334:19]
  assign topModule_io_inputs_3 = io_inputs_3; // @[TopModule.scala 370:23]
  assign topModule_io_inputs_2 = io_inputs_2; // @[TopModule.scala 370:23]
  assign topModule_io_inputs_1 = io_inputs_1; // @[TopModule.scala 370:23]
  assign topModule_io_inputs_0 = io_inputs_0; // @[TopModule.scala 370:23]
endmodule
